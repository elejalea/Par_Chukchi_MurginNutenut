Эвын И’УЛӃУТ
Лыги, лыгъоравэтльа ынкъаам айванальыт гэкрычмэ эймэвык, вама мэгчервагыргыт.
Ынӈин, ӄорагынрэтыльыт ӈэргэрык гавылгыӄаанмата, гырокы0ым гэкилвэе.
Айванальэн ынкъам лыгъоравэтльэн-аӈӄальэн гатвата Ръэвин крычмын – Полъа.
Ынӄэн, кэлик «Крычмыт айванальэн» Тасян Теин нивӄин, энмэн ынӄэн крычмын ынанъыттъыёл гамголен тааароӈо лыӈык айванальа.
Ынӄэн крычмын гэвытрэтлин унмытэленъеп рырынгээвынво ынкъам коргаво рытэ йитйив, пыкитльэн аӈӄальэты.
Чукоткакэн ынкъам Беринговкэн аӈӄак йитйив нывытрэтӄин гырокы ынкъам ӈэргэрык.
Ынкы наӈӄалӄатӄэнат аӈӄагыннэгӈыттыльыт.
Ыныкит ныръэвуӄинэт, ӄол нитӄинэт нъытвъэмэтӄинэт гаетъевма нымнымэты ныкэрэтъылёӈэт.
Наӄам ӄол ы’твъэт нынэквэтэвӄинэт аӈӄальэты ынпыначгынтанво, микынэ рырынгээвъёлӄыл рэмкыльын – йитйив кылетэ ымыльо таароӈвагыргыт аӈӄальэн.
Ынкатагнэпы нымгоӄэн крычмын Полъа.
