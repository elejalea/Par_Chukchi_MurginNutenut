Светлана КОЧНЕВА, заместитель директорэн Анадыркэн публичныкэн библиотекэн нынныльын Тан-Богоразын
Перевод Вама Майӈымараквыргын чукоткальыт гэпытлиӈичьэтэтлинэт тайкыма рэӈъатвывакъонвыт яанво ривлык риӈъэтвыт СШАйпы Советкэн Союзэты. 
Рэӈъатвыткоръэт Аляска –Сибирь гэтэйкылин 10 йъилгыӈит. 
Рэӈъатвывакъонвыт гамголенат тэйкык ымыльо ръэтык риӈъэтвыткукин. 
Нэкэм кытвагыргыт гэвытрэтлинэт Чукоткак, миӈкы тэӈвытку гамголенат тэйкык рэӈъатвывакъонвыт.
Нымытвальа Вэлӄылкин, Анадыркэн, Марковокэн, Чаплинокэн, миӈкы гатайкымголенат рэӈъатвывакъонвыт, ныйпэӄинэт рыпкэратъёттэ яанаӈат тарэӈъатвывакъонвыӈкэн ынкъам тараӈкэн. 
Нытъэрылтэтӄинэт мигчитльэт рабочийтэ ынкъам тарэӈъатвывакъонвыӈкы нывинрэтӄинэт ымыльо нымытвальыт, колхозникыт, служащит, рыбочийтэ, кэлиткульыт. 
Яанаӈат ныривлыӄинэт маглята.
Нэнакэтъатӄэн эрым эйгысӄыкин риӈэлейвыкин ръэткэн Герой Советкэн Союзэн Илья Павлович Мазурук: «Ынӈатал рэӈъатвыляйвыръэт Вэлӄыл-Красноярск колё нитчьэв гатвален. Ныриӈэмъетӄинэт лётчикыт чьэчеӈнутэйикви, энымкыльин, магнитныкэн компастэ ынкы мачьаӄаяаӈ нынъэлӄинэт. Плепы вальыт нутэкэлит лёӈытвальыт…»
Мачымыльо риӈъэтвык уйӈэ гатваленат энаномаваткэнат яанаӈат ынкъам рэӈаляйвыгыргын нымкыӄин лиӈыткучьывытгырӈит нитӄин гыйивӄэву катголтатгыргык лётчикэн. 
Маравыплыткок ынӄэн рэӈъатвыляйвыръэт гитлин тэнмычьо яамгок рэӈъатвыляйвыгыргын ынӄэн ныркывӄэн нутэйиквик.
Справка «КС»
Ӈыроӄ гивиӈит, октябртагнэпы 1942 гивикин октябртагнэты 1945 гивикин риӈъэтвыткульэ 1-ӄав Челгызнамяльын авиадивизиен гэныпкирэтлинэт АлСибъеквэ 8094 америкальэн риӈъэтвыт. 
Рэӈъатвырэвлыма гантымӈэвленат 81 риӈъэтвыт. 
Гараквачаленат 115 о’равэтльат.
