Гантэнмавлен Иван О’МРУВЪЕНА
Кэлиныгйивэтыльын Полина Александровна Максимкина гэпкитлин Чукоткагты 1933 гивик 18-ча элеӈитыльу.
Ынӈытэӄ редакциягты гатаписьмоӈлен ынинн ӈээкык Наталья Зорина, нымытвальын Хабаровскик, микынэ гатвыленат ытля ынкъам ытлыгын, мигчирэтыльыт ынкъам нымытвальыт Чукоткак гивиткуӈит, титэ тэӈвытку тъарваратыргэн нынтомгавӄэн калечетгыргын, титэ тэӈвытку гакалеткомголенат ы’ттъыютльэт игыркинэт эвынӈуткэкин нымытвальэн – винрэтэ русильин кэлиныгйивэтыльэ.
ПАЛЯНО НЪЭЙӇЭВӃИН КМИӇЭ
Наталья Зорина нытаписьм оӈӄэн: «Пыкиринэӈу Чукоткагты гымнин ытля Полина Александровна нивӄин, энмэн ытлён гамголен мигчирэтык ӄол чавчывэн нымнымык, вальын Увэлек чымче.
Ынкы нъэлык ынан янор нинэрэчичевӈиӄин нымытвальыт лыгъоравэтльат, наӄам люнрэӄыльэтыльын, аромкыльатка нытваӄэн, – нивӄин ыммэмы.– Кмиӈык ынкъам ыргинэт йытоткольык рээн тэрыгӈэ нымытвак, моонэн гыюлетык лыгъоравэтльэн йилыйил.
Йытоткольыт ивнинэт, иӈӄун вэлер ыннэн-ӈирэӄ лиӈыткучьывытгырык ыргынан ы’нытрилыркынэт кмиӈыт омакатынвы ӄол лыгэрак».
Янор калеткогыргын вэтгаво люӈылгыльын.
Авынчукоткальыт ынкъам ныӈинӄин кэлиныгйивэтыльын ӈэвысӄэтӄэй янор ыргичгу ныльувылгычичев вылгыӄинэт, ныйгулетӄинэт лыгъоравэтльэн ынкъам русильин йилымил яанаӈат.
Кэлиныгйивэтыльын кмиӈэ нъэйӈэвӄин Палейно.
1933-1934 гивиткуӈит ыммэмэнэ гыюленнин лыгъоравэтльэн вэтгав, кмиӈэ-ым – русильин.
1935 гивик ытлён нъэйӈэвын Анадырэты кэлиныгйивэтыльин конференциянвэты, ынӄоры нанъялгытатын нымнымэты Увэлен, миӈкы ынан льунин ы’вэӄучилӄыл Фёдор Зорин.
Чеэкэй моогъат кэлиныгйивэтык, Максимкина – лыгъоравэтльаелык.
Ӈинкэлиныгйивэтыльыт гэмигчирэтлинэт ымы Ӄытрык, нымнымык Пээк, ынӄоры Анадырык.
Еп пенсияльо энъэлкэ, Максимкина гитлин директоро Базовокэн калеткорак Анадырык, миӈкы нымигчирыйгулетӄинэт студентыт Анадыркэн педучилищакэн .
Мынивмык,1930-ӄав гивиткук Чукоткагты гэпкитлинэт ымы ӈавъелтэ Ольшевскаянтэ – Елена Фадеевна ынкъам Вера Фадеевна.
Ытри нэмыӄэй гэмигчирэтлинэт калеткораткок Чукоткакэн, Елена Фадеевна кэлиныгйивэтыльу, Вера Фадеевна – бибиотекак.
Чукотка ыргынан лёӈпэлята нэнтыгъэн, ӈутку гэпэлӄэтлинэт.
Пенсияльо нъэлык, Полина Александровна ы’вэӄучик ынкъам ытлювъёӄакйык рээн гаялгытлен Хабаровскэты.
Полина Александровна гаӈавытлювъёӄая нынымытваӄэнат ӈэранкомнатальын ярак.
Ыргин гатвален огород, миӈкы нынынӈэвӄинэт овощит.
Ныглёӄэнат Чукоткагты.
Нырэенӈыӄинэт титэ ӈан Чукоткагты.
Кытъаткэ-ым льэлеӈкы 2004 гивик ытлён уйӈэ нъэлгъи».
НЫМЫТВАВАГЫРГЫГЪЕТ ӇЭВМИРГИН
Рымагтэты Наталья Фёдоровна письмок гивлин: «Пээкик гым гъурэтигым 1939 гивик.
1946 гивик ытлыгын гакалеткомголен Хабаролвскыкэн парткалеткорак, кэлиткуплыткук ынкы гэмигчирэтлин инструкторо Крайкомык партиен, 1949 гивик-ым гэнӈивылин Чукоткакэн окружкомэты партиен, посёлкагты Анадырь.
Ыммэмы-ым, ӄонпы лымӈэнак мургин ытлыгык, гэмигчирэтлин кэлиныгйивэтыльу калеткораткок округэн.
Ӈавытлювъёӄай гымнин йытоткольэн Аня гэкэлиткуплыткулин пединститутык, гэнъэтлин кэлиныгйивэтыльу англияльэн ынкъам японыльэн йилык.
Ытлён энмэч ӈыроча гатвален Австралияк, Мальтак ынкъам Суматрак.
Ынӄэнат государствок ынан гэпирилинэт дипломтэ.
Ытлён мигчирэтыркын Хабаровскыкэн калеткорак.
Лыгэн-ым, ынан кылеркынин нымытвавагыргын ӈэвмиргин ынкъам мури мытэргавыркын.
