Светлана КОЧНЕВА, заместитель директорэн Анадыркэн публичныкэн библиотекэн нынныльын Тан-Богоразын
Ытлён гамэгчерымголен Чукоткак, титэ гэпкирлин 1955 гивик 18-ча элеӈитыльын.
Ӈотӄо ытлён Армиятванвэты гэпирилин.
Гэмигчирэтлин ывинтэтыльу ывэнтатрак, ымы рабочийыно, лымӈэ инженеро приискак «Отрожный».
Игорь Риган гатвален 23 элеӈитти, титэ ытлён гатвылен округкэн газетак «Советская Чуколтка»: «Акалырокыльэн, пэнин калевэтгавыльын, мытлётыльын, ӄэтпы корреспондент – ынӈин вальын ытлён.
Калевэтгавыльа лыги Игорь Рига – журналист округкэн газетэн.
Ыныкит ратвантык Эквыкыннотык, вэты ӄыйгулетгыткы ытлён.
Ынин варкыт тэӈкэлит, ымы ытлён таӈпычвэтгавтомгын, наранчаёвӈытык тэӈэвын».
Еп армиятвама ынан нинэнӈивыӄинэт калеёттэ вагыргыт маравратыльэн газетагты.
Декабртагнэпы 1959 гивик ынан моонэнат тэйкык материалтэ калейпатынво газетак «Советская Чукотка», ынӄоры гэкэлиткулин партийныкэн эквычьыкалеткорак отделенияк «Журналистика».
1971 гивик Игорь Рига гэнъэтлин члено Союзэн журналистэн.
Ынинэт тайкыёттэ вагыргыт гакалейпатленат газетак «Правда», «Труд», «Известия», «Комсомольская правда», «Магаданская правда», «Магаданский комсомолец», «Советская Чукотка», «Крайний Север», журналык «Политическая агитация», «Мир Севера», альманахык «Чукотка».
1976 гэвэтагнэпы Игорь Рига гамэгчерымголен Чукоткакэн округкэн нутэйгулеткин музейык.
Ынан гыёлятъёттэ вагыргыт вэты пэгчиӈу нылгыӄинэт ынкъам ныкалейпатӄэнат лымывнкы.
Ытлён гитлин редакторо икутъэр кэлик калеткольэты округкэн.
1981 гивик Магаданкэн такнигаӈынвык гэтэйкылин кэликэл Игорь Риган «Анадырь: историко-краеведческий очерк».
1990 гивик ынан гатвылен нымкыче вэтгавъёлгэпы «Анадырь – столица Чукотки».
Ытлён гэмигчирэтлин ымы телевиденияк, 2003-2004 гивиткуӈит нымкыче гатвылен ынӄо «История Чукотки глазами Игоря Риги».
2004 гивик ытлён гэнъэтлин дипломанто литературныкэн конкурсэн нынныльын Юрий Рытгэвын номинацияк «Докуменитальные истории», 2008 гивик-ым – эналватыльо конкурсык номинацияк «Публицистика» тэйкык кэликэл «Анадырь знакомый и незнакомый».
Ы’ттъыёлкэн часть кэликин гэтэйкылин Москвак 2009 гивик нъэлык 120 гивиӈитти столицэн Чукоткакэн.
Ӈирэӄэв часть кэликин ынан люӈыплыткутэ рыннин – ынӈингивик ытлён гэпэлӄэтлин.
Справка «КС»
Игорь Григорьевич Рига гинэнпиривлин диплома ынкъам знака «Лауреат премиен Чукоткакэн автономныкэн округгэн».
Ынин нынны гэкэлилин Анъякалек Чукоткакэн автономныкэн округэн, гинэнпиривлин лымӈэ знака «За преданность городу».
