Иван ОʼМРУВЪЕ
Перевод Хабаровскыкэн такнигаӈынвык «Гранд Экспресс» гэтэйкылин стихыльын кэликэл «Нас вдаль вела Полярная звезда».
Ынӄэн энмэч ӈирэӄэв кэликэл, миӈкы калейпатгъат стихыт эйгысӄыльин.
Ыʼттъыёлкэн ынӈин вальын кэликэл, миӈкы гатвыленат эвынӈуткэкыльин поэтэн тайкыёттэ, гэвытрэтлин 2017 гивик.
Ӈотӄэн туркэлик гакалейпатленат тайкыёттэ русильыйиле тастихӈыльа, нымытвальа Чукоткак мэчынӈытэӄ.
Наӄам русильин поэттэ этлы ытръэч нытастихӈынат, лымӈэ ытри нитӄинэт йилыльэтыльу эвынӈуткэкыльин тэкэлиӈыльин – лыгъоравэтльэн, айванальэн ынкъам ӄаарамкэн елепы.
Ӄымэлым калевэтгавыльа, нымытвальа Чукоткак лыги нэтчынэт эвыӈуткэкыльин поэттэ.
Йилыльэтыльу итыркын ымы Андрей Носков, микынэ гэнумэкэвлинэт тайкынво кэлик стихыт эвынӈуткэкыльин.
Ынан гэйилыльэтлинэт русильыйилымил тайкыёттэ лыгъоравэтльарык Пётр Оʼмрынтона, Вера Иʼвӈэвытынэ, Валентина Иʼтэвтэгнынэ (Вэӄэтынэ), Александр Аʼтавӄайына ынкъам Елена Оʼмрыӈана, ӄаарамка Андрей Кривошапкинына ынкъам юкагирыльа Николай Куриловына.
Тывъёлӄыл, пэгчиӈу таӈылгыӈ тайкыёттэ кэлик магаданыльа Сергей Сущанскийына, микынэ нымкыӄин гивиткуӈит румэкэвыркынинэт вагыргыт тэкэлиӈыльин Северо-Востокэн Россиен.
Ынӄэнат нэмыӄэй гакалейпатленат туркэлик.
Ӄымэл-ым игыркин калевэтгавыльа лыги рэтчыгнин, ынӈатал кытвагыргыльо гитлин калейпатынвы ыргинэт тайкыёттэ вагыргыт.
Лымӈэ кэлик гакалейпатлен повесть туртэкэлиӈыльин «Оленные люди» («Чавчыват») Вера Грачёван.
Поэзия туркэлик рывэнтыркынин вальа Майӈымаравынвык поэта Борис Боринына (Блантер), мэӈин горатвален мигчирэтык редакцияк округкэн газетэн.
Юрий Рытгэвынэ, Альберт Мифтахутдиновына ынкъам Виктор Кэвылӄутынэ рээн гэргыпатленат туркэлик поэттэ Михаил Эдидович, Анатолий Пчёлкин, Татьяна Ачиргина, Илья Юрьев (Логинов), Геннадий Сабанцев, Олег Комаренко ынкъам ӄутти, микынти лыги нэлгыркынэт мурыгнутэк ынкъам микыргин тайкыёттэ ӄол гитэ кытоор гакалейпатленат округкэн газетак «Крайний Север».
