Иван ОМРУВЬЕ
«Лыгъоравэтльат ынӈатал пэнинэт мытлёчетовэчватыльыт, – кэлик гивлин эргыпатыльын учёный Владимир Тан-Богораз. 
– Галяк ӈроӄ– ӈраӄ ы’лёӈэттэ эмнуӈкы лымэвыр аӈӄачормыкэ ытри нъирэӄинэт, гэнпэ амалваӈ вальыт рыпъёт и’гнэлгыт, нэннэтнэлгыт ымы. 
Лымӈэ ытри гарачвыӈа, гэтэйкэвэ, гэпиӈкучитэ ынкъам ӄутти». 
Мытлёчсетовэчвыт гэкэлилинэт 1979 гивик тэкэлиӈыльэ Владилен Леонтьевына кэдлик «Ынанкатгочьын, ынанмылычьын».
Чаата гинэкынъучитэ. 
Ӈаргын гумэкэтэ ӈинӄэгти ынкъам гамгота увичвэтык. 
Нытвэтчаӄэнат эмтъэръюну ӈирэӄ амъянра увичвэтыльыт ягна ыргичгу, ыргин вытгыргыпы ӄол увичвэтыльын рынныа’мата гакынгынтыгалята, ӄол гитэ гэнвилысӄычетэ лымэвыр ынан гэтиӈусӄычетэ а’матъё рыннытъол, ныппылюӄин отгэты акынъокэгты. 
Ӄутыргин чааттэ кытчымча нирӄинэт айъока а’матъё рыннылгын, элвэльинэргин-ым ынраӄ гэнармагта а’матъёк. 
Ынанэнакынъочьыт гакоргава инэкынъук. 
Ынӄэн увичвэт нытвыӄэн ӄорачет. 
Гымнан тыкэтъоркынат увичвэттти ӈинӄэю вамакэн. 
Энмэч мытлыӈгэвэльо ынпыянва нынинъэйвымури гырыткук, ымыльо гачаата ӈинӄэйин. 
Пууръу рынык ӄулин гъэмэтэ, гэрэкынъуӈэ выроттыӄагтэ, мэчемгитлеӈин. 
Ӄулин пууръу увичву гэлгэ рырамавъё тэвъэл. 
Микынэ нинэкынъуӄин, ынӄэнына нинэнуӄин тэвъэлытъул.
