Светлана КОЧНЕВА, заместитель директорэн Публичныкэн библиотекэн нынныльын Тан-Богоразын городкэн Анадырь
15 июнык эвынӈуткэкыльин поэтэн, тамэнӈымлявыльэн ынкъам актёрэн Виктор А’рэчайвынэн (1937-1993) 80 гивиӈитти о’раттагнэпы.
Виктор А’рэчайвын гъурэтлин Эӄӄэник, вальын аӈӄачормык чымче Льорайпы (Чукоткакэн район). 
Ынан гэкэлиткуплыткулин Анадыркэн педагогическыкэн училище Айгысӄываратыргэн, миӈкы эӈъэлю рытчынэн тэӈыйгулетык поэзия ынкъам млявыт ченэтваратэн. 
Кэлиткутумгык рээн ынан нинэтэйкыӄин журнал «Юность». 
1957 гивик тэминӈычьэтыльын студент лыги рытчынин эргыпатыльа дальневостоккэн поэта ынкъам йилыльэтыльэ Валентин Португаловына. 
Ытлён нэмыӄэй гантэнмавлен акватынво чукоткакэнат ӈиныльык рээн VI Ымнотаеквэкэн фестивалеты ӈиныльин, э’митлён гатвален Москвак 60 гивиӈитти яалегты – 1957 гивик. 
Ынӄэн ӈиныльин крычмынвык А’рэчайвынына рыкалыровнэн чиниткин мляв «Собачья упряжка» ынкъам «Фестивальная песня», э’митлён ынӄоры гэйилыльэтлин Валентин Португаловына, калейпатъё ӄутти кэлик ынкъам чукоткакэн литературак. 
Фестиваль рыгъевавынво А’рэчайвынына гантомгавлен ӈирэӄэв мляв «Трубка мира».
Кэлиткуплыткук педучилищек А’рэчапйвын ганватлен Аӄӄанэгты, гитлин заведующино нымнымкин клубык. 
Ынӈингивиткук ынан моонэнат кэлик лымӈылтэ. 
Ынӈот гивлин кэлиныгйивэтыльын Льурэкин калеткоракэн Изабелла Автонова: «Талпыӈӈок 1960-ӄавкэнат гивиӈитти нымным Эӄӄэни гатвылен пэлянво нымытвальа, ынкэкинэт о’равэтльат ганъялгытавленат Льорагты. 
Виктор А’рэчайвын ӄитпэквъи ынкы нъэлык рытомгавынво грапчакэн-млявкэн ансамбль Аӄӄанэльэпы. 
1969 гивик коллектив гантомгавлен нымнымкин Льурэкин Ярак культурэн. 
Ансамбль говэчвынкалыровлен Анадырык, Магаданык, Москвак, гатвален Аляскак (США). 
Вараткэн коллективо гэтэныннынлин 1975 гивик».
Грэпыт ынкъам млявыт, тайкыёттэ Виктор А’рэчайвынына 1970-1980 гивиткуӈит ынкъам рыкалыровъёттэ лыги гэтчылин ымыльы Чукоткаеквэ. 
Чывипыт грэпин «О новой жизни» гаяален овэчвынкалыровкэн программак Государственныкэн лыгъоравэтльэн-айванальэн ансамбля «Эргыръон».
А’рэчайвынына лыги гэлгылин онмэргыпатыльын тамэнӈымлявыльын Нутэтэгын, мэӈин нэмыӄэй гатвален VI Ымнотаеквэкеэн фестивалык ӈиныльин ынкъам студентэн, нымикыче ыныгрээн говэчвынкалыровлен.
Виктор А’рэчайвын лымӈэ эргыпатыркын ӄнур актёр, мэӈин гувичвэтлин ӈыраӄ художественныкэн кинофильмык: «Начальник Чукотки» (1966), «Самые красивые корабли» (1972), «Кит и компания» (ГДР, Чехословакия, СССР, 1974) «Смок и Малыш» (1975). 
А’рэчайвын гитлин магляльо ынкъам винрэтыльу эргыпатыльэты америкальэн грапчальэн ынкъам актёрэн Дин Ридына кинок «Кит и компания», тайкыё кэлигйит Джек Лондонын. 
Кино тайкыма гаяален ы’ттъыгаканъе А’рэчайвынэн.
Виктор А’рэчайвын гэпэлӄэтлин 1993 гивик, 56 элеӈитыльу.
