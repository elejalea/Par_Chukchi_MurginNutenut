Дина КЭУКЭЙ, авынбиблиограф анадыркэн Публичныкэн библиотекэн нынныльын Тан-Богоразын
Амрытэнма 20 сентябрык  1648 гивик ыʼтвэ Дежнёвын гагалялен Майӈыэʼӈыткын.
Ынӈингивик русильин аӈӄаляйвыльа гэмо гэлгылин, иӈӄун гатвален эргыпатыльын м айӈывагыргын – гэныгйивэтлин вальын  иʼрвытгыр Евразиен ынкъвам Америкэн.
Мытлыӈэн гивиӈитти галягъат, титэ 26 сентябрыу 2013 гивик экспедиция «Арктика– нутэйиквин гыюлеткин» гэпкитлин Анадырык, эʼмитлён гатвылен газетак «КС».
Ынӈингивик ӈирэӄ уттъытвэ «Святитель Николай» ынкъам «Апостол Андрей» наяагъан аӈӄаляйвыръэт, тэӈвытку яаё Семён Дежнёвына Тиксэпы Анадыртагнэты.
Тэнмычьын «Арктика – нутэйиквин гыюлеткин», рыкытвылявъё эмвинрэтык Русильин географическыкэн обществота ынкъам Правительствота Чукоткакэн, пэгчиӈу гэлгылин общественностя ынкъам гитлин гыёлятъёно кытвагыргыт российскыкэн Арктикэн, гэнанкэтъоӈатлен эргыпатыльык вагыргык российскыкэн историен ынкъам географиен, гинэнӄитпэвыткулин раройвавынвы вэнратвылгыгыргыт ыргичгу регионтэ экономическыкэн, научныкэн, культурныкэн ынкъам тунриистическыкэн вагыргык.
Мынынкэтъоӈатын, элек 1648 гивик ыннанмытлыӈэн ыʼтвыт, миӈкы гаӈатваленат вальыт экспедицияк Семён Дежнёвын ынкъам Федот Поповын тэӈвытку гэлейвылинэт Чукоткакэн аӈӄаеквэ, микырык нагалянат амрытэнма ыннэн тысяча километртэ аӈӄагычормыеквэ.
Гыёлятъё вагыргыгъет, Беринговкэн эʼрвытгыртагнэты гэпкитлинэт ӈыроӄ ыʼтвыт, ыннэн гэпылӄэтлин иʼрвытгырык.
Энмэч Беринговкэн аӈӄак ӈэргэрык эйичгэ ганъянръавленат гынульыт ӈирэӄ ыʼтвыт.
Поповын ыʼтвъэт гагчорматлен вытгырык нотачьомыткынтэ Дежнёвын ынкъам Чукоткакэн танкавӈынво чимэтыльын ыʼтвъэт ынкъам мимлыйырэтык аймыёчгыт.
Эвынӈуткэкыльык рээн маравпэнрыткок ытлён гатынвылен.
Дежнёв ынкъам ынинэт 25 лейвытумгыт ганомленат Олюторскыкэн нотачьомыткынык.
Галяк вытку 10 неделят аӈӄаляйвыльыт гэпкитлинэт Анадырык.
Семён Дежнёв ынкъам 17 казакыт гэльэлеӈитлинэт 1648-1649 гивик Анадырык, миӈкы нэтэйкынэт еп эръилекэ вээм ыʼтвыт.
Элек 1650 гивик, тылек гыргочагты Анадырваамэн пыльыльыайгыпы наянат ыргынан 600 километртэ.
Ынӈэнӄач Дежнёвына рытомгавнэн льэляӈэтваны, ӈотӄоры тывъё Анадыркэн острого, русильин авынванво Чукоткак XVII-XVIII столетияк.
Семён Дежнёвына гэтэйкылин нутэкэликэл Анадырваамъёчгэн (гантымӈэвлен).
Элек 1652 гивик Анадырваампыкэргырыкэн нотачьомыткынык гэльулин рыркаровтын.
Элек 1660 гивик пууръу Дежнёвына эрму гэнъэтлин элвэльин оʼравэтльан, ытлён-ым тумгык рээн гаваӈӄынма нутэйиквитэ чейвэ гэквэтлин Аколымагты.
Аӈӄаляйвыльа Семён Дежнёвына ынкъам Федот Поповына, ыргинэт лейвытумгырык ганръачӈытовлен ымнотаеквэкэн эргыпвагыргын: нэныгйивэтын иʼрвытгыр Азиен ынкъам Америкэн, нэнвэнтын Северо-Востоккэн нотачьомыткынык Чукотка ынкъам нанъомравын ынӄэн нотачьомыткын Русильин государствэн Тихий аӈӄачормык.
Лымнʼэ
Галяк 120 гивиӈитти, 1898 гивик, ванляк Русильин географическыкэн общество, ынаннэкъаяӈӄачкэн нотачьомыткын Азиен гэныннэтлин «нотачьомыткыно Дежнёвын».
