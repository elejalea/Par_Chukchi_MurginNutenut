Гантэнмавлен Вадим НИКОЛАЕВЫНА
Перевод Лыгъоравэтльэн, о´птыма ӄнур ӄолеваратэн, нэмыӄэй гатвален эӄунмэтйильыт нэмык´эй нытэнымчеӈӄинэт.
Ынӄэн вагыргын ыргынан кытэ нынръачӈытовӄэн, титэ алваӈ а´анляӈ.
Ӄол ынӈин вальын вагыргын гатваален ынкъам гэкэлилин 1955 гивик, ганымӈылявлен нымытвальа Нунъэмук Константин Иивынэ., э´митлён гавалёмлен ынан  ынпыянвэпы аӈӄачормыкэн Беринговкэн и´рвытгыркин.
Вагыргын гакалейпватлен номерык 1 «Записки Чукотского краеведческого музея», тайкыё Магаданкэн такнигаӈынвык 1958 гивик.
Ынӄэн гатвален лыгитэленъеп.
Пинакулык, Ӄытрык ӄача, гэльэлеӈитлин америкальэн шхуна Ынӈингивик лыгъоравэтльаваратэн гатваленат ытръэч пойгыт ынкъам ырытти.
Шхунак-ым гатваленат мушкетти – милгэрти.
Шхунак гэмигчирэтлин матросо –ӈуутвыльу лыгъоравэтльан-чавчыв.
Ӈэнку ытлён нанмыгъан.
Гэетлинэт чыченткинэльыт тымъён, ыргынан намӈылёнат ы´твыльыт.
Капитана гочленат:
– Гэмо, миӈкри ӄытгъи.
Йъилгын галягъэ, ӄол лыгъоравэтльата гэлкытлин, мэӈин тэгинӈэтыльу гитлин: ӄол матроса мынга рыкалыровнэн тэгинӈэтыльын капитан, рыгивэннин, миӈкри тымъё лыгъоравэтльан мэмлыткынэты гэнинтылин.
Ынӄэн лыги лынъё вагыргын-тагэнӈатгыргын ганымӈылявлен ӄотырыкы томгэты-лыгъоравэтльэты.
Гыттэпычьын нутэтумгын гивлин:
– Рэ´итыгъэ аӈке´ы, ытри ралвавӈыт ӈотӄо ы´твыткук.
Моргынан мытранмыӈын капитан, амыргынан матростэ мытранпэлявӈынат.
Ыргынан нанмыгъан ыннэн о´равэтльан, ымы морнынан мытранмыӈын ыннэнчьэн.
Инъэ капитан охотанвэты ӄытгъи.
Ынкы лыгэн варат ӄутгъи натваалынат ырытти гамъамэма.
Лыгъоравэтльа нэйпыгъэн тыляръэт капитанэн ынкъам ӄолентогъат.
Гыттэпычьын гивлин:
– Ӄырыткутык ынӈэн мачогты, ипэ нанӄэты, ӄэлюӄ тымнэн ынапн рэӄык лёӈэнаачьыльын, тымӈэтвальын.
Лыгъоравэтльат ырыткугъэт.
Капитан ыннанванвык вакъогъэ, люӈӄулильэтыльын, ипэ гинрынин мъамэлгын атынвэпы.
Ынкы лыгъоравэтльарык ынкъам пойга нанмыгъан.
Капитан нэнумкэвын лыгъоравэтльамэл., нэвиръытвыгъэн ынкъам эвиръыт ынан яаёттэ олёвынвык нэтрилынэт.Эргатык лыгъоравэтльа найъогъан ы´твъэт ынкъам ӄолентогъат:
– Ӄыйъогыткы чиниткин капитан ынкъам ӄыгитэгыткы.
Моргынан ытлён мытынмыгъан, мури эмэлкэ гэӄунмэтйимури.
Ынкъам ы´твъэт эквэтгъи.
