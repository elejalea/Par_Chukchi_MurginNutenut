Иван О’МРУВЪЕ
Перевод Мытлын’эн гивин’итти галягъат, титэ 17 январык 2013 гивик ганъомравлен Постановление правительствэн РФ рытомгавынво национальныкэн парк «Берингия».
Ынк’эн пууръу чит вальын региональныкэн паркык ынкъам нъэлгъи федеральныкэн парко.
К’ол ынкэкин участокык, еп антомгавка парк, гым гатвайгым 60-к’ав гивиткук XX векэн.
Ынк’эн Чагтоваамъёлгык, ипэ-ым Чагтоваампыкэргыргык, мин’кы гатвален нымным ан’к’агыннэгн’ыттыльэн.
Нымнымык чымче вээмк’эйык к’ача гатвален пограничникын застава, мин’кы гым нъармиятвайгым.
Оттырак’айык нымнымкин нынымытвак’энат колхозникыт.
Мургин заставак гэтэйкылинэт казарма, элгытавран, тылячьыран ынкъам к’утти имыръэкинэт оттырак’агтэ.
Ваамк’аеты наймыморэ, мин’кы э’лк’эпы нэнакаймэморэ э’лен’н’эк’эгти.
Ынн’ингивик гым люнчимгъульигым, ынк’эн рэк’ыннык’эгти мыткаймэркынат.
Амынан ныкоргавморэ льук ынк’энат э’лен’н’эт.
Элек-ым Чегтувээмык йин’э ныкин’вин’умури, ынн’атал нычачак’энат.
Мимыл-ым вээмин нычык’к’ин ынкъам эн’уйкыльин, о’птыма лелелк’эргычьыпэральын.
Гымнан ымы игыр, галяк нымкык’ин гивин’итти, тытан’кэтъоркын ынк’эн ваны, Чегтувээм пыкирыльын Чукоткакэн ан’к’агты.
Этааны, тымн’ъатав лён’ынтымлявыльын Чагтоваамъёлгын паркагты «Берингия», э’митлён вэты тан’ыйголятъёлк’ыл ынкъам гытамо лынъёлк’ыл.
Справка «КС»
Ымыльэты нутэйиквин паркэн 1.819.454 гектармэл кывальын.
Паркык варкыт мытлын’эн лымынкы вальыт участоктэ, нак’ам амчекыяа нымнымыткойпы нутэйиквик н’ырок’ муниципалитетэн Чукоткакэн АО.
«Колючинский», «Чегитунский», «Дежнёвский», «Мечигменский» ынкъам «Провиденский» – гамгаучасток ыннаны апэракыльэн.
Паркагты гантымлятленат илирти: Аракамчечьын, мин’кы варкын ровтын рыркэн ынкъам гылмэмлыванвыт; Ы’ттъыгран – ынкы варкын «Китовая аллея», рытомгавъё амрытэнма мытлын’эн вектэ яалегты; ваамъёлгын Чегтукин – гыргоча ынк’эн вэмин гэльутэ кытэпат: илирти Литке ынкъам Беннета, кынман’к’ы Лаврентия ынкъам к’утти ванвыт, э’митлёнат вэты тан’ыйголятъёлк’ылтэ.
