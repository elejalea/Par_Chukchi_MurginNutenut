Иван О’МРУВЪЕ
Перевод Лина Тиӈыл гъурэтлин ройыръкык ӄорагынрэтыльэн. 
Гэкэлиткуплыткулин 1956 гивик Ленинградкэн педагогическыкэн институтык нынныльын Герценын. 
Гитлин воспитателё калеткорак илиркин Аён, лымӈэ кэлиныгйивэтыльу Анадыркэн педагогическыкэн училищек Айгысӄываратыргэн. 
Январык 1970 гивик Тиӈыл гэльулин председателё исполкомэн Чукоткакэн округкэн Советэгн депутатэн мэгчетльываратэн. 
Гэӄитпыльэтлин Лина Григорьевна рытаӈытватынво вэлыткогыргын ынкъам о’рамръагъепыткогыргын ӄорагынрэтыльык. 
Сессиянвык масӄонпыӈ вэтгаво нылгыӄин энантаӈытватгыргын национальныкэн нымнымыткук. 
Лиина Тиӈыл ынкъам ӄутти члентэ исполкомэн нытгымэтӄинэт, иӈӄун тараӈыльа вэты лыги ы’нылгыркынэт эвынӈуткэкинэт ӈаргынэнавагыргыт тараӈма. 
Гэӄитпыльэтлин винрэтык поэто нъэлык Антонина Кымъытваал.
1983 гивик Магаданык гатвален Ымроссиякэн семинар ӈиныльин литераторэн Эйгысӄыкин, Сибиркэн ынкъам Дальний Востоккэн, миӈкы вэтгаво гэлгылин ымы гымнин тайкыё повесть. 
Ынӈингивик Лина Тиӈыл нымигчирэтӄин лыгъоравэтльаелымэл редакцияк Магаданкэн такнигаӈынвыкэн ынкъам гэӄитпыльэтлин семинарынвык. 
Ынкы вэтгаво гэлгылин ымы гымнан калеё вагыргын колхозаткэн. 
Лина Григорьевна гивлин: «Ӈотӄэн кэлик плепы тывыркыт ымыльо вагыргыт чавчывэн, мургинэт ӄорагынрэтыльэн. Колхозатгыргын кэлик еп микынэ нымкъэв атвыка ынкъам пагчеӈгыргын, иӈӄун О’мрувъена мэчтэӈвытку ынӄэн кэлинин. Ӄэлюӄ-ым ытлён вэты мыкмигчирэтыльылӄыл тэкэлиӈкы, гыюлетыльылӄыл…».
