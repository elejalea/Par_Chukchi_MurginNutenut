Вера ТЭВЛЯНТО, урэмигчирэтыльын қорагынрэтгыргык, Эквыыннот
Перевод Талпыӈӈок февральининик март эмнуӈыльыт нытэнмавӄэнат Тэркыӄаматынвэты, ыьтри ныялгытӄэнат торавээнвэты, торралӄаӈынвык нытаароӈӄэнат, ялгытыркыт торавээнвэты, торралӄаӈынвык таароӈыркыт, рагролмын гытамо нэлгыркын миӈкриым эргатык рэмкын льаляӈэтынвэты ратэнмавӈыт.
Еп рэювкы вулӄытвик ӈавэтынва етьа рытчыркынин рэнтыткоолӄылтэ нотатаароӈкэн льаляӈэтынвэты.
Ройыръэн эвиръыт рытэнмавыркынэнат, инъэ таӈгаглыйпы.
Етьа рытчыркынинэт уттыт увинтэткин ынкъам гытамэты рытрилыркынинэт этролклыӄылтэ.
Ы’ттьыт омрыквотыркынэнат аръасэнтыкэгты.
Ӄэлёӄ-ым гытамо нылгыӄинэт, нэкэм таароӈыӈӈок.
гыгэру ныльгыӄинэт ымы мэйӈыӄулильэтык. Ынкъам нывириӈкинэт майӈывэтгавыльыт.
Кимылтэтыльыт экэвку нылгыӄинэт, нэкэм ӈэвъэнйыръыт.
Инъэ ривыльэ рыпкирэтыркынин ӈэлвыл, лыгэнэвыт ӄутти ӄлявылтэ гырыткугилиркыт.
Эвыт тангиянъё кынъоёлӄыл ӄораӈы эвытрыкэ вак, э’ми ӄаачыкогты ныргэлӄин, - лыгэнэвыт ӈавэтын нъэйӈэльэтӄин.
Ръэнут винвынъэӄэрэвын, иа’м тыӈэво лыӈыркын, эвытлым винвъутык титэ.
Ыныкит пэлле аймэтъёлӄыл ныкынъуӄин, ынпыначгыт ныринӈычьэтӄинэт.
Ымылыгэн аманъята нытчыӄин.
Тиркыӄэмэтык ачгыта чама тымӈалголяӄ ныръилеӄинэт.
Нутрии ымӄэтпыльата нитӄинэт ымы ынпыначгыт, ымы мыӄыльыт.
Майӈыӄылявылтэ ныгагчавӄэнат корагыркэнвэты, ръэлятэнмавыркыт.
Чымӄык а’ачегъянвыт рачвыӈыркыт, пэӈкорачвыӈыркыт.
Тэӈычьу нылгыӄин элёльычетгыргын.
Ӈутку ымы мыӄыльыт гэчевкы нытваӄэнат нэкэм эпэрык рээн.
Чьэчеӈкы нывириӈӄинэт рыровэты рачвыӈыльыт, энмэн рыӄывэтоӈыт, аӈъачгыргын вээнток.
Мыгрэмкыльэтык гэчевкы рэмкын ныльувылгыӄинэт.
Ынпыначгыт, ынпыӈэвэ гэтэнгиеӈэ ӈэвычӄэтти ынкам эккэт гэныгивэтэ.
Нээккэльыт-ым гарыглята - вэчьым ӈээккэт нэтэныггивӈыркынэт.
Энмэч-ым ӄутти гаӈавынрагтата.
Лымӈэ
Тэеӈкы янот – ым ялгытыӈок ынпыначгыт чимгъуркыт,парыркыт, нэныгивэвыркын льаляӈэтынвылӄылтэ.
Элгулеӄ-ым лымэвыт ильуткуркын, эвыт вак ярартамэнӈыльын.
Ыргынан нэльуркынэт лымкэты вальыт ванвыт льаляӈэтынвыкэн.
