Иван О´МРУВЪЕ, пограничнико гитлин
Перевод Пириплыткук город Кёнигсберг 1945 гивик 33-ӄав мотострелкакэн полк маравратыльэн НКВД гэргыпаныннатлен «Кёнигсбергский».
Энмэч маравыплыткокэнат гивиткуӈит Кёнигсбергскыкэн орденыльын Красной Звезды пограничникэн отряд ганъялгытатлен Чукоткагты, э´митлёнын штаб гатвален нымнымык Гуврэл (Урелики) Провидениякэн районкэн.
Пограничникэн армиятвагыргын гатвылен журналистарык, маравратыльа, историка ынкъам ымы Игорь Ригана.
Э´квыргъам игыр мытытвыркын энакэтъатгыргын вагыргыгъет армиятвакэн ынӄэн эргыпатыльын пограничникэн отрядык.
Ӄутти нутэтумгыт гъармиятваленат ынӄэн пограничныкэн отрядык, ымы рыпкэратъёттэ мэйӈынутэкин нымнымыткойпы, микыргин ытлыгин ынкъам миргин энъататгыргын маравынвык гатвылен журналиста, тэкэлиӈыльэ, лымӈэ кэлик историкын ынкъам краеведын Игорь Риган «Анадырь знакомый и незнакомый».
Кытоор гым нэмыӄэй гъармиятвайгым ынӄэн пограничникэн отрядык, гатвайгым мачымыльо ан+ӄачормыкэнат нымнымыткукин заставак, ымы вальын э´ӈыткынык Халюскиын.
Игыр ынӄэн застава уйӈэ, ымы ӄутти чит вальыт.
Игыр армиятвальэты пограничникэты винрэтыльу нутэгынрырэтык итыркыт технологическыкэнат яанаӈат, пограничникыт-ым чит вытэчгыргыпэральыт эвиръыльыт паагъат армиятвак нымкыӄин нымнымыткук, миӈкы кытоор гатваленат застават.
Э´ӈыткынык Халюскиын гынрырэткин ваны гатвален энмыткынык, миӈкы гырокы ынкъам ымаляӈэт галегӈытота амалваӈ вальыт галгат, Армияплыткоӈӈольыт нылиггичиӄинэт ынӄэнат рырагтатынво майӈнотагты.
Тыкэтъоркын, Халюскинкэн э´ӈыткынкэн заставак гъармиятваленат сержант Галацан, старшина Родионов, рядовойтэ Батурин, Зуев, ынӈин нынныльын эрым заставакэн старший лейтенант Зуев.
Гымнан лыги, ыргинэт ытлыгыт, миргыт, йичьэмиттумгыт, чакэттыт гатваленат Майӈымаравынвык вэрэӈынво чычетнутэнут пэнрыткольэпы а´ӄальэпы.
Лёӈынтыяата тынтыркынэт ымы нутэтумгыт ыӈэн отрядык армиятвальыт: сержант Николай Макотрик, рядовойтэ Виктор Татыга, Николай Тэвлянто, Иван Никулин, Александр Гэматагын ынкъам Иосиф И´нмугье, ефрейтор Сергей Кымъылгын,..
Лыги тылгыркын ымы ваӈӄыттамэнӈыьын, эргыпатыльын художник Россиен Иван Сейгутэгын, мэӈин нэмыӄэй ӈроӄ гивиӈитти гъармиятвален ынӄэн пограничникэн отрядык.
Галяк нымкыӄин гивиӈитти, энмэч армияплыткотагнэпы, титэ нытэнмавэгым 2001 гивик риӈэк Франциягты, таӈавэтываӄ тыльугъэн ӄлявол, мэӈин нэмыӄэй гъармиятвален заставак, вальын э´ӈыткынык Халюскинын.
Горатваморэ пычвэтгавык, гакоргавморэ, оптыма чычеткинэльымури!
Гым гъармиятвайгым ымы заствак вальын нымнымык Чегтун.
Ынӈэнӄач аркын вээм, ынӈатал чыӄмимлыльын, мэйӈылыгинныльын, ӄнур гытгыткок Ватыркакэн эмнуӈкы, миӈкы ымы варкыт кычавыт, туйкэт, ӈэгныкин-ым вээмыт лымӈэ гаварэӈочьыленат.
Чегтук нытумгыльэтигым ӄутти нымытвальык рээн.
Гымнан а´ӄантыяатыӈ армиятвагыргын Кёнигсбергыкэн пограничникэн отрядык, э´митлён гантомгавлен 75 гивиӈитти яалегты, титэ гамаравпэрэлен мурыкэкыльэ город Кёнигсберг.
Справка «КС»
20 сентябрык 1945 гивик комиссра НКВД СССР гэнынныкэлилин приказ рытомгавынво 33-ӄав ӄэгнэвыткукин полкэпы Кёнигсбергыкэн орденыльын Красная Звезда пограничникэн отряд, э´митлёнына гынрыру лынъёлӄыл нотачьомыткын Чукоткакэн.
26 отрядык 1946 гивик штаба отрядэн, вальын Провиденияк, заставальэты ынкъам ынкъам комендатурэты приказ гынрырэткин нотачьомыткынык.
Горатваленат вак оьтрядык 21 застават, миӈкы гатваленат ынкы армиятвальыт о´равэ\тльат.
Ынӄоры ынӄэнат рытъэрытвэвэ гэнтылинэт.
1967 гивик пууръу комендатурак гэтчылинэт группат, заставак-ым эмрынгиитэ гамголенат гынрыру лыӈык.
Ынкатагнэпы гамголенат гынрыру яау тылячьыяанаӈат вэтгавъёлгыльыт.
1990 гивик Анадырык гантомгавлен комендатура, миӈкы гатваленат ӈирэӄ застават.
2005 гивик гаялгытатлен ымыльэты отряд Анадырэты.
Игыр ынкы армиятваркыт пограничникыт, микырык эмӄынгивик 28 маяк нэкрымыркын Ы´лёӈэт пограничникэн, титэ вэты наэргыпавыркынат ыргын ы´ттъыётльат о´равэтльат.
