Григорий ТЫӇАНӃЭРГАВ, нотагаймычьыэнарэрыльын
Перевод Гымнан лыги тылгыркын, ръэнут нытвыӄэн гымнинэт йытоткольа Эналватык э´ӄэльык. 
Ынӄэн гымнан а´ӄантыяатыӈ, миӈкри ӄун ытлыгын ынкъам ытля ынӈатал гакытрэватленат вэнратынво нутэвмрмӈэтыльыт. 
Гымнан тыкэтъоркын, иӈӄун ынпыянвыт, ӈинӄэю нъэлык гачечавыӈӈойгым, ӄонпы кытрэвчемгъогты нытваӄэнат валёмтагнэты, титэ мурыгнутэльэ налвын фашизм (нотапэнрыткольа э´ӄэльыт). 
Йытоткольыт ынкъам чычеткинэльыт нонмыкытрэватӄэнат мигчирэтык, ыргынан ымы гым гынрыру люӈылгэ: ынанъыттъыёл гэчимгъутэ рымкэвык ӄаат, ӈаргыночьыналгыт мыкыӈ рытчык, ныкэрэтъылёӈэт тэйкык лилит, кълит, эвиръыт, плекыт. 
Ынӄоры ымыльо тайкыё миӈкриӈан нынэквэтэвӄин (нивӄинэт, энмэн нотавэрэӈатыльэты), иӈун пытӄымгок ванӈэлтатык.
Ынӄоры кытваӈэлтатык паагъат ымыльо, нивӄинэт, мараквыргын паагъэ, мурыкэкыотыт эналватгъат. 
Ымы гым коргыӈ тынъэлык. 
Ытлыгын ынкъам ытльа гинэнпиривлинэт гомударственныкеэн медаля Амэналватык э´ӄэльык.
