Дина КЭУКЭЙ, авынбиблиограф анадыркэн Публичныкэн библиотекэн нынныльын Тан-Богоразын
Кэлиныгйивэтыльин, журналистэн, поэтессан Тамара Кликунован (литературныкэн пытӄынынны Смолина. – Прим. ред.) 7 июлык нъэлгъэт 80 элеӈитти.
Ялгыык Анадырэты ыʼвэӄучик рээн, Кликуновырык эӈэлю гэлгылинэт рыкытвылек икутъэр райъонъёлӄылтэ кмиӈырык. Ыргынан ымваӈэт ӄитпу гэлгылин  кмиӈин литературныкэн-публицистыкэн студия «Умка-пресс» ынкъам гэтэйкылин гыюлеткин кмиӈин журнал «Умка», китӈин литературныкэн журнал «Муракашка», лымӈэ икутъэр сборникыт кмиӈин.
Кликуновынтэ  инъэтэтык 1992 гэвэтагнэпы округкэн эвыннымнымык эӈъэлю гэлгылинэт рылек Ыʼлёӈэттэ славянскыкэн письменностэн ынкъам культурэн.
Ынанъыттъыёлкэн кэликэл Тамара Кликунован «Лунный иней» гэтэйкылин Анадырык 1996 гивик.
Галяк-ым ӈыраӄ гивиӈитти Москвакэн такнигаӈынвык «Магазин искусств» кынмал Владимир Кликуновына рээн гэтэйкылин кэликэл «Подарок Полюса Надежды».
2005 гивик Тамара Кликунова гэнъэтлин дипломанто гыёлчетгыргык «За образцовое владение русским языком в профессиональной деятельности» мэгчетльэты кэлиныйгулевкин Россиякэн Федерациен, 2006 гивик гаянотлен журналистэн конкурсык «Отражение», 2010 ынкъам 2014 гивиткук нъэлгъи дипломанто литературныкэн конкурсык нынныльын Юрий Рытгэвын.
2010 гивик нъэлгъъи члено Союзэн писателен Россиен.
2009 гивик Новосибирскыкэн такнигаӈынвык гэтэйкылин ынин кэликэл «Карусель» курэ чиниткин манэта.
Галяк ӈыраӄ гивиӈитти Москвакэн такнигаӈынвык «Спутник» гэтэйкылин кэликэл «Мне есть что вспомнить», миӈкы гатваленат стихыт ынкъам пыӈылтэлтэ.
Ынӄэн кэлик гакалейпатленат эргыпатыльыт Чукоткак оʼравэтльат Маргарита Глухих, Валентина Вэӄэт, Зоя Ненлюмкина, Михаил Меринов ынкъам ӄутти.
Чымӄык вагыргыт калеткоракэн гатвыленат разделык «Дневник учителя».
Разделык «Из блокнота журналиста» гатвыленат  таӈъоравэтльат Чуоткакэн.
2015 гивик Новосибирскыкэн такнигаӈынвык «Гео» гэтэйкылин кэликэл «Тропинки к юности», миӈкы гатваленат 23 рассказтэ.
Кэлиныгйивэтыльын, журналист, ӄэтпъоравэтльан – ынӈатал наройвыӄэн ынӄэн ӈэвысӄэт, пэнин тэӈычьэтыльын  нымытватомгэты, ымыльорыкы.
Ымы игыр, энмэч пенсияльо нъэлык, лёнтымӈэтвата итыркын, ӄонпы ринъэтэнӈыркын имырэӄык.
Справка «КС» Тамара Николаевна Кликунова – лауреат премиен Магаданкэн комсомолен, Тэминнʼыльын вараткэн кэлиныйгулевкин,  урэмигчитльэн Россиен, урэмигчитльэн Чукоткакэн, гинэнпиривлин Анъякалета Думэн Чукоткакэн АО.
2007 гивик Тамара ынкъам Владимир Кликуновынтэ гинэнпиривлинэт ордена нынныльын князыргэн Пётр ынкъам Феврония Муромскийыргэн кʼитпинъэтэтыльыт мигчирык ынкъам энанъомравыльыт ройыръынымытвак.
Майык 2015 гивик Тамара Кликунова гинэнпиривлин энакэтъаткэн гиивкʼэвэ рырынгээвма 85 гивинʼитти оʼраттагнэпы Юрий Рытгэв.
