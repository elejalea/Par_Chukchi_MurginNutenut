Дина КЭУКЭЙ, Иван О´МРУВЪЕ
Перевод Моотагнэпы Ы´ттъыёлкэн Камчаткакэн ляйвыгыргын Витус Берингын ынкъам Алексей Чириковын 24 январык рэнъэлӈыт 295 гивиӈитти (1725), гыму лынъё ынкъам рывъёльавъё Петербургыпы Пётр Великийына гыёлятнво ванвыт, миӈкы Азия «гатымлятлен Америкак ынкъам мэӈӄо таӈыпкэрыӈ городэты европальэн».
Ынӄэн ляйвыгыргык Ы´ттъыёлкэн Камчаткакэн эрму гитлин датчаныльын Витус Беринг, мэӈин еп 1704 гивик гаялгытлен Россиягты.
Мурыгнутэк ытлён гэргыпатлен гыютльу аӈӄаляйвыльо петровкэн флотэн.
Ляйвынвык ымы гатвален онмэргыпатыльын гыютльэн Алексей Чириков.
Ляйвыма ынан гэкэлилинэт вагыргыт лейвыкин.
Учёныйырык гэйгулетлин аӈӄачормыеквэн Майӈыгэляӈӄэн, гэнумэкэвлинэт ынкъам гэйгулетлинэт ӄутти вагыргыт эвынӈуткэкыльин, нымытвальэн Эйгысӄынутэк ынкъам Дальний Востокык, гэвилыткупууръыткулинэт варатык рээн ынкэкин, лымӈэ лыги гэтчылинэт ӄутти вагыргыт вилыткукин Америкак ынкъам Японияк рээн, ӈаргынэнакэнат вагыргыт гэйгулетлинэт, Эйгысӄыкинэт гынникыт, гэкэлилинэт вагыргыт Востокэн Сибирэн, лыги гэтчылинэт ляйвыръэттэ ӄутти нымытванвыткогты, вальыт чекыяа.
Галяк вытку ӈирэӄ гивиӈитти ляйвыгыргыльыт гэпкирлинэт Охотскык.
Вытку июлык 1728 гивик ы´твъэт «Святой Гавриил» гаӈӄалӄатлен райъоӈынво и´рвытгыр Азиен ынкъам Америкэн, гатваленат лейвыльыт кынмаӈӄак Креста, бухтак Преображения, нэнвэнтын илир Святого Лаврентия, ынӄоры натагъан и´рвытгыр, э´митлён ӈотӄоры гатвыӈӈолен нынныльу Берингын.
Лейвыльэ гэтэйкылин аӈӄакалекал, миӈкы гатвыленат льоёттэ нотачьомыткынтэ Чукоткакэн, Кагынинын, Чаплинын ынкъам ӄутти.
Нутэкэлик лымӈэ ганкалыровлен, энмэн Чукоткакэн нутэнут миӈкы лёнтымлятыльын.
