Гульнара СИБГАТУЛЛИНА
Талпыӈӈок январь Ассоциациен эвынӈуткэкыльин нъэлгъэт 28 гивиӈитти рытомгавтагнэпы.
Ынӈингивиткуӈит ынкэкинэт членыт ынкъам ӄитпыльыт гинъэтэтлинэт рыплепавынвы нымкыӄин вагыргыт нымытвальэн округык.
Ассоциация имырэӄык гыюлетгъи ынӄэнат ӄымэк 30 гивиӈинӈит.
Ымы эргыпатыӈӈогъат, ӄэтпымэгчерыӈӈогъат общественныкэн вагыргык ӈиныльыт.
Саша Тэвлявъе игыр итыркын ы’ттъыёлкэн вице-президенто Ассоциациен, мэӈин еп энма студенто эвын гэӄитпэвлин инъэтэтык общественныкэн мигчирык.
- Тэӈвытку гым общественнико гитигым еп 2002 гивик вэрэӈынво правот ынкъам вагыргыт айгысӄываратыргэн, титэ гэкэлиткуйгым Санкт-Петербургык.
Ынӈингивиткук Ассоциацията тъарваратыргэн нинэнумэкэвӄинэт ӈиныльыт ванво семинарык,миӈкы нинэйгуленмури вагыргыт мургинэт, тъарваратыргэн, - нивӄин ытлён.
- 2005 гивик, титэ гатвайгым Анадырык, нымкыӄин вагыргыт тытэӈыйгулетынэт, ынӈингивик гитигым винрэтыльу Управлениягты КМНЧ Аппаратэн Губернаторэн ынкъам Правительствэн Чукоткакэн АО рылянво Совет выёльыргэн авынчукоткальэн.
2007 гивик Александра гэнъэтлин члено президиумэн, гитлин секретаро, 2011 гэвэтагнэпы нъэлгъи члено, инэнлельу ӈиныльин вагыргык.
Ынӈингивиткук ӄитпыльыт, миӈкы гатваленат Виктория Анака, Анатолий Ӄэргынват ынкъам ӄутти – ныӄитпыльэтӄинэт рылек эмыръавагыргыт ӈиныльин: курсыт гыюлеткин чычеткин йилык, крычмыт, мытлёчетгыргыт, ӈаргынэнагынрыраткэнат общественныкэнат мигчитти.
Игыр авынтэнмычьо мигчирык Ассоциациен итыркын «Школа молодого лидера», э’митлёнын 2017 гивик нъэлгъэт мытлыӈэн гивиӈитти.
Ынӈингивиткуӈит мыкыӈ 150-к ӈиныльыт ым-Чукоткакэн гинъэтэтлинэт ынкы.
- 2015 гэвэтагнэпы гымнин общественныкэн мигчир мыкэтгъи.
Игыр эӈъэлю мытылгыркынэт вэрэӈъёлӄылтэ правот эвынӈуткэкыльин кылек ымыльо вагыргыгъет ыргинэт, - гивлин рымагтэты Александра.- Яачыӈкэнат 5-7 гивиӈинӈит мургин Ассоциацията эӈъэлю рытчынинэт нымкыӄин мигчитлыӄылти, э’митлёнат ӄутти энмэчевын пэгчиӈу ынкъам инъэтичгу нэтчынэт – ынӄэн «Э’раӄор» ынкъам «Э’йӈэв».
Наӄам ӄоргаво мытылгыркын, иӈӄун ынкы гиливыркыт мыкыӈ эвынӈуткэкыльыт, нымытвальыт нымнымыткук мурыгнутин.
Вице-президент лымӈэ гивлин, иӈӄун игыр Ассоциацията тэӈынчичьэтыркынин нотаяакэн вопрос.
Ынӄэн чимгъуу лыӈыркыт ынныӈыттыкинэт участоктэ, гыннигӈыттыкинэт, лыгэн-ым нотаяакэнат вагыргыт.
- Мургинэт райъонъёлӄылтэ пэнинэт.
Коргаво мытылгыркынэт о’равэтльат, организацият , винрэтыльывт Ассоциациягты рэнъатытвэвынво ымыльо вагыргыт эвынӈуткэкыльин, - плытковачык гивлин Александра Тэвлявъе.
Справка «КС»
Ассоциация авынчукоткальэн гантомгавлен 28 январык 1990 гивик.
Чукоткакэн АО ынӈингивик гатымлытвален Магаданкэн областэты.
Ы’ттъыёлкэн эрму ынкы гитлин Александр О’мрыпкир.
