Светлана КОЧНЕВА, такалгын директорэн Анадыркэн публичныкэн библиотекэн нынныльын Тан-Богоразын
15 гивиӈитти галягъат (2002), титэ Увэлек гамголен тэйкык ынаннэкъаяӈӄачкэн православныкэн часовня (таароӈран). 
Увэлен варкын нивлыӄин тэпӄэк, Чукоткакэн аӈӄачормык. 
Сентябрык 2002 гивик ынкы гамголен тэйкык православныкэн часовня (таароӈран) Воскресения Христовын.
Гэнанмыгоӈатлен тэйкык таароӈран-кэтъоран Губернатор Чукоткакэн АО Роман Абрамович. 
Тараӈыльо гитлин тараӈкэн предприятие Омскэпы. 
Таароӈран гэтэйкыплыткулин 2003 гивик.
Тывъёлӄывлтэ ӈирэӄ ынӈингивик вытрэтыльыт вагыргыт. 
Ынӄэн гэльулин этлы амтараӈыльа, ымы Увэлельэ, микырык мычвыно натчыӈӈогъан таароӈатгыргын. 
Титэ намгон тэйкык яраӈы, люур вай айгысӄыӈӄач вытрэтгъи тиркыӄымчучьын. 
Ганоратвавлен эмилетык рыгырголявык крест гонпыма. 
Титэ-ым мигчир нэплыткун, таӈавэтываӄ тэӈмэлетгъи ӈаргынэн. 
Ынпыянвыт нивӄинэт, ынӈин тэӈвытку вагъэ, миӈкри ӄун ипэ нъэӄэйгэтыркын. 
Лыгэн-ым вагыргыт ынӄэнат ӄэглынангэт гатваленат.
