Гантэнмавлен Дина КЭУКЭЙЫНЭ, Иван О´МРУВЪЕНА
Перевод Ӄол ынанъыттъыёлкэн гыю- летыльин Сибирык Семён Дежнёвын ӈутингивик нъынъэлынэт 415 гивиӈитти о´раттагнэпы (1605–1673).
Айгысӄы-нэкъаяӈӄачкэн нотачьомыткынык Чукоткакэн гэтэйнылин кэтъоквын ынӄэн эргыпатыльэн ноталяйвыльэты–аӈӄаляйвыльэты Рэӄэ гэргыпатлен Семён Деэжнёв, ръавагырга – ынкэгйит пыӈылтэлыркын москвакэн тэкэлиӈыльын айгысӄывагыргыгъет Вячеслав Огрызко.
Гъурэтлин Семён Дежнёв нымнымык Осиновская Двинскыкэн уездыкэн ройыръык аӈкальэн, – гэкэлилин ынан. – 25 элеӈитыльу гатвален Тобольскик.
Яачы гэнӈивылин Енисейскэты.
Эйгысӄынутэк тэӈвытку гатвален 1638 гивик, титэ отрядык рээн казакэн Посника Иванова Губаря гатвален ноталяйвынвык Янагты ынкъам Индигиркагты.
Дежнёвына гэльулинэт амалваӈ вальыт ынкъам нымкыӄин вагыргыт ноталяйвыма.
Нымкыче ытлён гапэнрылен Вытку ытлён гатынлен 1641 гивик.
Ынӈингивик Дежнёвына ынкъам ӈроӄ казакырык рээн рыльатэнма налог Якутскэты.
Ынӄэн пэнрыма ыныкы ытлён ӈирэче гатынлен.
Ынӄоры гатвален ляйвыгыргын Оймаконэты, миӈкы нэмэ ытлён ганроӄавлен атынык.
Еп атвака Оймаконык ынан гэльулин якутӈав Сичко Абкаяда, микынэ гагтолен ыныкы экык Любим.
1643 гивик Дежнёв Михаил Стадухинына рээн гэлейвылин пыкэргыргыпы Алазеян пыкэргыпгытагнэты Экулымэвээмин, миӈкы нэтэйкын льэлеӈиткин нымным, э´митлён ӈотӄоры ганъялгытатлен ваампыкэргыгэты Сухой Анюй Акулымагты.
Ынӈин гатомгатлен нымным Нижнеколымский, э´митлён гэнъэтлин авынбазано ӈотӄокэнат экспедицияльэты, мэӈо нымгоӄэнат налогэнарэркэнат ляйвыгыргыт.
Кытъаткэым льэлеӈкы нэмэ гатвален ынин кытвагыргын.
Нымнымэты гапэнрытколенат мыкыӈ 500-к юкагирыльыт.
Дежнёв гатынлен левтык мъэмитэ.
1648 гивик Дежнёв ытри Федот Алексеев Попов тэӈвытку гаталенат кочаы´твэ э´рвытгыргыпы Азиен ынкъам Америкэн.
Кытъаткэ а´нӄагыргын ляйвыгыргын вама гатвален этчывагыргын: эйичгэ лымынкыри ганлыплятленат ы´твыт казакыргэн.
Ӈыпэльыт Дежнёв ынкъам икутъэр казакыльыт аӈӄачормык вытку январык 1649 гивик чейвэ гитлинэт пыкэргыргэты Анадырьваамэн.
Льэлеӈитыльыт, титэ гэквэтлинэт 13 о´равэтльат, нэтэйкын коч-ы´твъэт, рэӄэ гырголятгъа ваамъеквэ гырголятгъат, миӈкы натайкымгогъан ӄол нымным, э´митлён ынӄоры гатвыӈӈолен Марковоно.
Вээмчурмык Анадырь Дежнёв гатвален 12 гивиӈитти,миӈкэкин варат налогпэрэёно гэтчылин, ынкэкинэт лыгъоравэтльат.
Ӈотӄоры ынан тайкымгоёттэ нымнымгыпы гэквэтлинэт экспедицият К. Ивагновын Х 1660 гивик кынмаӈк(´агты Крестэн, ынкъам кынмаӈӄагты ПровиденияЪ Л. Морозкон ынкъам И. Голыгинын (1685 гивик э´ӈыткынэты Олюторский) ынкъам В Атласовын (1697 гивик Камчаткагты).
Рымагтэты Вячеслав Огрызко нымӈылтэлӄэн, энмэн 1662 гивик Дежнёв ганватлен Якутскэты, ынӄо ытлён нэнэквэтэвын Москвагты.
Столицатагнэты ытлён гэлелин мыкыӈ ӈирэӄ гивиӈинӈит.
Москвак гаманэмынгыквын ытлён 19 гивитуӈит нутэлейвыкин ынкъам аӈӄаляйвыкэн: 28 рублти, 22 алтынтэ ынкъам 39 манэт, лымӈэ 97 аршинтэ сукнота.
Ынӈин гаймычьыпэрэк Дежнёв ынӄоры нэмэ гэквэтлин Якутскэты, миӈкы гэӈирэӄэвлин ӈавтыӈык амынан нъалыльэты чит ӈэвъэнин пылвынтытамэнӈыльэн Арбутовын – Кантеминкагты Архипована, микынэ гагтолен ыныкы экык Афанасий.
1666–1668 гивиткуӈит Дежнёв гэмигчирэтлин вээмык Оленёк.
Ынӄэн ваампыкэргыргыргын гэльулин тэӈвытку еп 1620 гивиткук Иван Ребровына.
Янор ынӄэн микырык пэгчиӈу люӈылгыльын.
Чекалваӈ пэраӈӈогъэ вагыргын, титэ ваамэты Анабар пыкиргъэт мангазейскыкэн казактэ.
Сибирскыкэн властя гэтчылин ӈэранчывэӈ Анабарскыкэн-Оленёкскыкэн район.
Тунгустэ, вальыт чымче гытгык Ессей, нагынрэтыӈӈонат Магазеяльа, оленёкскыкэнат-ым тунгустэ – Якутыльа.
Воеводтэ Мангазейкэн ынкъам Якутскыкэн ӄонпыӈ нынмаравчеткэнат ыргичгу, иӈӄун ытри таӈналогпэрэӈ.
Амынан Дежнёв гэтъивыльэтлин вагыргыт маравчеткэн амаравчеткэнано рытчык.
Тэнмычьо, ынан ганпааӈатлен чит вальылӄыл пэнрыткогыргын боягтарыргэн оленёкскыкэ тунгусэты.
Гэпэлӄэтлин Дежнёв 1673 гивик Москвак.
Справка «КС»
Энмэч 1736 гивик Г. Ф. Миллеоына ынанъыттыёл сибирскыкэн архивык гэльулинэт челобитныйыт (калеёттэ вагыргыт).
1910 гивик яатльарык мурыгнутэкин э´ӈыткынык нангырголявын рэргыпавынво русильин аӈӄальын уттэ тайкыё крест.
