Василий И’УЛӃУТ
Перевод Таӈоонъынтаӈ нъэлгъи. 
Мыкуунъыльын мургин эмнуӈ. 
Оонъыгэчегыргын нэмыӄэй гыму гэлгэ эвынӈуткэкыльэ, иӈӄун ынӄэнат рук ымы льэлеӈкы. 
«КС» калейпатыркынэнат икутъэр тэтлегмимлыӈкин тэнмычьыт оонъэпы калейпы Изабелла Автонован «Авынроолӄылтэ лыгъоравэтльэн ынкъам айванальэн».
ЭТЛЕГМИМЫЛ РЫВАРЭВЫЧЬЫЛГАВ ЫНКЪАМ РЫСАХАРЭЛГАВ
5 кг вэривычьин, 1 кг сахарэн, 1 чаёкэн вонны гвоздикэн, 10 л мимлин. 
Ымыльо ынӄэн чыӄмэмлыттъыёлӄыл, энааръёлӄыл сахара, гвоздиката ынкъам а’тчаёлӄыл 19 ы’лёӈэттэ, этлегмимыл таӈылпыӈ нъэли.
ЭТЛЕГМИМЫЛ РЫВАРЭВЫЧЬЫЛГАВ
150 г уунъин, 120 г сахарэн, 1 л мимлин. 
Ынӄэн етъаӈ рытчыё пъэттыёлӄыл. 
Ынӄоры гылмэмлыттъыёлӄыл ынкъам рэтэтъёлӄыл 5 мин. 
Уунъыт ититыльыт атлягмэмлепы рыъянръавъёлӄылтэ. 
Этлегмимыл рыӄытвэвъёлӄыл. 
Таӈылпыӈ ынӄэн галяк 1-2 ы’лёӈэттэ.
ЭТЛЕГМИМЫЛ РЫВАРЭВЫЧЬЫЛГАВ ЫНКЪАМ РЫМЁДЫЛГАВ
150 г вэривычьин, 150 г мёдэн, 1 л мимлин.
Рытэнмавык тэкэм энмэч ы’ттъыёл тывъёмэл, ытръэч пууръу сахарык яаёлӄыл тэтлегмимлыӈык мёд.
ЭТЛЕГМИМЫЛ «УТРО»
1 стакан этлегмимлин рыварэвычьылгав, 1 чаёкэн вонны кофеен, 1 чаёкэн вонны сахарэн. 
Ынӄэн рэтэтъёлӄыл ынкъам аӄытвэкэгты пыльёлӄыл.
