Светлана КОЧНЕВА заместитель директорэн Анадыркэн публичныкэн библиотекэн нынныльын Тан-Богоразын
85 гивиӈитти галягъат, титэ 24 мартак 1933 гивик ганъомравлен мэгчертэнмычьын Челгыракэн.
ЫМГЭВ ЭӇЭТ ЛЕЙВЫЛЬЫН ЛЫМЫНӃО
Культбазат гантомгавленат вэнратынво аӈӄальыварат Чукоткакэн.
Чавчыват-ым вэнратынво III съездык Советэн Чукоткакэн районкэн 1932 гивик гавэтгыльатленат делегаттэ ванляк Дальневосточныкэн Комитет Эйгысӄин ынкъам Чукоткакэн окрисполком мачалваӈ рытчык культбаза, иӈӄун чымчаӈ нымытвальык, ымы чавчывак рытчык ынӄэн.
Ынӄэната 24 мартак 1933 гивик гантэнмавлен тэнмычьын рыялгытата рытыльын политикакэн-просветительныкэн учреждеие, тывъё Челгырано, эʼмитлён гиливыльылӄыл Ынаныяакэн Эйгысӄык.
Ынанъыттъыёлкэн Челгыран гэвытрэтлин Чукоткакэн культбазак рыкалейголявынво чавчыват, 1940-ӄавкэнат гэвэтагнэты Челгырат гантомгавленат ым-Чукоткаеквэ.
Челгырат гиливыльылӄылти ымгэвэӈэт, ялгытляйвык лымынӄо, эʼӄу рытчыёлӄылтэ ынӄэнырык эӈэӈыльыт, вэнратъёлӄылтэ ынӄэнырык ӈэвысӄэтти ӄитпэвык общественныкэн митгчирык, инъэтэтыльылӄылти рывантынво калеткорат ынкъам ынкы кытрэватыльылӄылтэ ымыльо нымытвальыт, рыкалейголявъёлӄылтэ ытри.
Калейголятгыргыт нынлеӄинэт чычетйиле – лыгъоравэтльэн, айванальэн, ӄаарамкэн, миӈкы ныйгулетӄинэт ванвыкэнат партиякэн мигчитльэт.
МАНЭНОМАКАКВЫРГЫН ЫНКЪАМ КУЛЬТУРАВАГЫРГЫТ
Майӈымараквыргын вама рывэтгыльаквыргыгъет крайкэнат комитетэн партиен гэнымкэвлинэт Челгырат, чит 1940 ынӄэнат гатваленат 24, 1944 гивик-ым энмэч 37.
Ынкы мигчитльэт мыкыӈ гэнъэтлинэт , кэлит гэнымкэвлинэт яанво.
Майӈымараквыргын вама Челгырат ынкъам изба-читальнят гинъэтэтлинэт ромакавынво манэт нотавэрэӈатыльэты.
Тэнмычьо, заведующина Челгыракэн Рыркайпиякэн сельсоветэн И.И.Рэнтыгыргына 60-ча гэнумэкэвлинэт нымытвапльыт тывынво Майӈымараквыргын, нотавэрэӈатгыргын.
Ынин бригада гатвален 14 нымнымыткук, ӄымэл-ым гэнумэкэвлинэт 2925 ӄорат нотавэрэӈатыльэты.
1949 гивик Рывэтгаквыргыгъет Советэн Министрыргин СССР законо гэтчылинэт челгыральыт вэнратынво ӄорагынрэтбригадат.
Челгыральо гэтчылинэт лымӈэ кэлиныгйивэтыльын-библиотекарь, фельдшер ынкъам киномеханик.
Мараквыргын плыткук Челгыральа тъиву гэтчылин нинъэйвыткумигчир нымытвальык.
Ынӄэнат гатгэлевыӈӈомголенат ӄорагынрэтбригадак ынкъам уткучьыткульин ванвык.
Челгыральа тъиву гэтчылин культурамэл энанпаӈъэвӈытоквыргын ӄорагынрэтыльык, ынныӈыттыльык, гыннигӈыттыльык, лыги лыӈык вытрэльыт ымнотаеквэк вагыргыт.
Нэкэм гэтэӈмигчирэтлинэт Нутэпынмыкин, Илирӈэйкин, Энмыльыкэн Челгырат.
Ынкэкинэт мигчитльэрык эмнуӈкы нынлеӄинэт экономикагъеткэнат семинартэ, ныныпкирэтӄинэт ӄорагынрэтыльэты газетат ынкъам журналтэ, нынпалёмэлявӄэнат эмнуӈыльыт вэтгавъёлгэпы вэтгавыльыт чычетйиле.
Чымӄык Челгыральа нытэйкыӄинэт газетат.
Заведующий Нутэпынмыкин Челгыракэн Нутэтэин гинэнпиривлин ордена Трудового Красного Знамени.
Справка «КС»
Культуракэн-гыюлеткин учрежденият Чукоткак гэнымкэвлинэт: 1952 гивик 75 учрежденияк культурэн гэмигчирэтлинэт 148 оʼравэтльат, ынкыгрээн 55 эвынӈуткэкыльыт.
Клубык, Челгырак, изба-читальняк гамэгчерымголенат гыютльэт оʼравэтльат.Майык-ноябрык 1949 гивик Анадырык гатваленат курсыт культурамэгчетльэн Челгыракэн.
Гэпкитлинэт Чукоткагты майӈынотайпы специалистат, Ам-1959 гивик Чукоткагты гэнӈивылинэт 32 гыютльэт культурамэгчетльат.
