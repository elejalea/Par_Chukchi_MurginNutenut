Светлана КОЧНЕВА, заместитель директорэн Анадыркэн публичныкэн библитотекэн нынныльын Тан-Богоразын.
14 июлык гэнъэтлинэт 95 гивиӈитти эвынӈуткэкыльин нымнымин Вэлӄыл Эквыкыннотыӈӄач вальэн. 
1922 гивик айванальа, нымытвальа Уназикык, гантомгавлен аӈӄачормык Крест нымным Вэлӄыл. 
Ӈотӄоры ырыкы чеэкэквъэт ӄутти ройыръыт нутэтумгин. 
Вэлӄылыльыт нымэмылӈыттыӄэнат, нырыркаӈыттыӄэнат, ныръэвӈыттыӄинэт. 
Ынкъам ныкимитъылпууръыткуӄинэт чавчывак. 
Советкэн вагыргынляма нымнымыльэ нынмэйӈэвӄинэт риӄукэт гыннэграк. 
Ныгынритӄинэт элгартэ, нымигчирэтӄин ваӈэран. 
Вама Майӈымараквыргын вэлӄылыльыт нэмыӄэй гакытрэватленат мигчирэтык вэнратынво нутэвириӈэтыльыт ынкъам лывынво э’ӄэльыт нотапэнрыткольыт.
Игыр Вэлӄыл эргыпатыркын, лыги нэлгыркын мургин нутэ-
тумгэ – вама Майӈымараквыргын ынкы гэтэйкылин рэӈъатвывакъонвын, мэӈӄо нынтакаӈатӄэнат Аляскайпы риӈъэтвыт тыляма рэӈаръэтъеквэ Аляска-Сибирь (АлСиб).
Маравыплыткокэн гивиткуӈит ынӄэн нымнымык гатваленат пограничникыт, олёвынвык гэтэйкылин кэтъоквын рэргыпавынво риӈъэтвыткульыт раквачальыт. 
Кэтъоквын игыр гынрыру, гытамо нэлгыркын Вэлӄылкин кэлиткульэ.
Вэлӄыл ык гэргыпатленат: Лейта-Тъаю – инэнлельын ансамблен «Имля»; Ким Акилькак – орденыльын Трудового Красного Знамени, ынанъыттъыёлкэн председатель колхозэн «Угляткак»; Василий Ятыргын – итыльын председателё сельсоветык, тэкэлиӈыльын; Михаил Ваалгыргын – аӈӄагыннэгӈыттыльын, член Союзэн писателен СССР.
Справка «КС» Нымным Вэлӄыл варкын 100 километрмэл урэльу посёлкайпы Эквыкыннот, айвачыӈӄач э’ӈыткынык Аннюалькаль кэтэм аӈӄачормык. 
Нымным гэтэнынныӈлин Вэлӄылю ванвык ръэвин вэлӄылмил пэральык.
