Григорий ТЫӇАНӃЭРГАВ, нотагаймычьыэнарэрыльын, г. Анадырь
Эргыпатыльа геолога Григорий Андреевич Тыӈанӄэргавына тывыркынэн кытооркэн чиниткин мэгчерымгогыргын геолого итык.
– Ынанъыттъыёлкэн гымнин нотагаймычьыэнарэргыргын гатвален ваамнолгык Алярмаут, айгысӄыӈӄач игыркин городык Билибино.
Ынӈингивик еп уйӈэ гатвален город.
Мури Сеймчангыпы мытинмык риӈъэтвэ Черскийтагнэты, вальын Экулымэк.
Ынӄо самолёта АН-2 мытинмык базатагнэты ГРП Каралваамкэн.
Ынкы гырокы гэмкэтлинэт отрядтэ аʼтчальыт рэӈанво мэгчерванвытагнэты.
Ымы мури.
Ӄынвэр нэмыӄэй мытриӈэмык.
Еп авакъока мытльун гырголяйпы вакъонвык рыгъеватъё крест, энмэн ӄырымэнаморэ вакъольылӄылморэ.
Ӄэлюӄ-ым мытынванмык, мэӈӄо ӈан гэриӈэмури.
Еп рэӈатыляма ӈэнри эрым отрядэн гивлин, чейвэ итыльылӄылмури базатагнэты.
Ынӄэн 100 километрмэл урэльын ръэт.
Лыгэн-ым мытимтинэт имтитэючгыт ынкъам мытэквэнмык чейвэ.
Ӈыроча мытыткивмык тылянвык.
Пыкиринэӈу мытымӈылёгъан эрым, иаʼм нанъотавмык вакъок.
Ытлён гачыӈытколен ынӈот: «Нъатчальатэгым, титэ рэпкиры самолёт, ыннээн-ым галяркын… Тынныӈыттымгогъак аʼтчама тури, Этъопэл гымыгрээн вакъок. Юрэӄ-ым алваӈ ратвагъа…».
«Ръэнут алваӈ нъытвагъан» – ынӄэн лёӈытва рыннин.
Геолого энма гым нымкче гитигым риӈъэтвэ, мачам-АН-2-а.
Риӈъэтвыткульыт гагтывэнратленат нотагаймычьыэнарэрыльэты нутэлейвык.
Наӄам ыргынан нынвакъовӄэнат риӈъэтвыт тымӈалголяӄ миӈкы, кытвыл атыроочгыкэванвык.
Лыги тылгыркын ынӈатал тэминӈыльын риӈъэтвыткук Борис Комков – нывэймэнӄин оʼравэтльэты, пэнин коргычьатыльын.
Ыныкит гырголяйпы эльукэ нинэнтыӄин кавэты вальын вакъон, етгыр нэнанвакъовӄэн АН-2, нивӄин, иӈӄун рымагтэты чейвэ мынинмык, гивэ морыкы: «Имтитэ рымагтэты ӄитгытык - акэмылтаткэгты мэгчерынвэты».
Ӄэглынангэт, ынӈатал ынан гэтэӈийгулетлин мигчир геологэн.
