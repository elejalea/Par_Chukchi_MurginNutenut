Иван ОʼМРУВЪЕ
Перевод Ынинэт тэӈкэлит такнигаӈынвык пэтле нытэйкыӄинэт 100 тысячтэ мыкэльу. 
Журналистэн, тэкэлиӈыльин Анатолий Ваховын 8 февралык нъынъэлынэт 100 элеӈитти оʼраттагнэпы (1918-1965)
Ынинэт кэлит мыгъянва чит пэнинэт калевэтгавъёттэ. 
Ымы гым ныпэгчиӈэтигым корынво ынӄэнат, ынӄэната вэлыткорак нынъэлигым, титэ нэнавалёмэгым, иӈӄун ынӄэн рывэлытковынво ганатвыленат кэлит, миӈкы гатвылен ыʼттъыёлкэн Ревком Чукоткакэн – «Ураган идёт с юга» ынкъам «Утренний бриз». 
Ыʼттъыёлкэн кэлик Ваховына плепы гатвыленат кытвагыргыт энантомгавкэн вараткэн вагыргынлягыргын ынаннэкъаяӈӄачкэн нутэйиквик Россиен. 
Ӈирэӄэв кэлик «Утренний бриз» рымагтэты гатвыленат ӄутти членыт ыʼттъыёлкэн Ревкомэн Чукоткакэн, советкэн оʼравэтльат энанаройвавыльыт нутэйиквик Ынаныяакэн Эйгысӄыкин. 
Вагыргыт гражданскыкэн маравмакэн гатвыленат ӄол кэлик Ваховына – «Адъютант».
Вахов гъурэтылин Дальний Востокык, ынӄэната мачымыльо кэлик, ынан тайкыёттэ, гатвылен ынӄэн нутэйиквин ынкъам ымы аӈӄы. 
Ӈинӄэйтумгык рээн ытлён нымкыче гэттэтлин ӈэйык Тигровая, мэӈӄо нытэӈвытрэтӄин Уссурийскыкэн кынмаӈӄы. 
Ӄол боцмана нэнатвыӄэнат аӈӄаляйвыгыргыт. 
Аӈӄы чимгъучыку гэтчылин ӈинӄэе. 
Боцман-ым ӈайгпы Тигровая гэкэлилин кэлик «Трагедия капитана Лигова» ынкъам ынкы гэныннэтлин Ходовыно.
Тэкэлиӈкы Вахов гамголен пэтле, ынинэт кэлиткукинэт сочиненият ынӈатал иничгыту ынкъам пэгчиӈу гэлгылинэт ӄутырык, калеёттэ мачалваӈ тэнмычьыкэнак тасочиненияӈкэн. 
Еп аʼачеко ытлён гэчимгъулин нъэлык журналисто.
Ынинэт кэлит, гэчевкы вальыт, нытэйкыӄинэт такнигаӈкэн ванвык нымкъэв. 
Ымы игыр ытлён накалевэтгавыркын, ӄэлюӄ ынинэт кэлик гатвыленат вальыт кытоор вагыргыт мургин дальневосточныкэн нутэк.
