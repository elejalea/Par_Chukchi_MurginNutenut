Ӄутти  эвынӈуткэкыльин лымӈылтэ игырыткукин калевэтгавэльа тымӈъатаво гарылга. 
Лыги лынъёлӄыл: ынӄэнат лымӈылтэ  кмэӈэты гатва, чама гэйилыльэтлиинэт росельыелепы гаглеты. 
Эʼквыргъам вэлер-ым ынӈин, ӄэлюӄ гатвыленат мургинэт ыʼттъытльэрык ынкъам варатэн гаймычьо итыркыт. 
Игыр ӄол лымӈыл мытытвыркын. 
Пипикылгын тымкыгэн'гыпы нылейвыкин. 
Пипи¬ӄылгэ льунинвэлвын, эйӈэвнин:
– Апай, ӄыетги, мымлюгыт!
Ӄытгъи вэлвын. 
Пипиӄылгэ мылёʼ'ӈонэн. 
Мылёма йылӄэтгъи вэлвын.
Лыгэн йылӄэтгъи вэлвын, льулӄыл кэлийвынин пипиӄылгэ вэлвын вылӄэ. 
Льулӄыл кэлийвыплыткунин, эквэтгъи пипиӄылгын. 
Йылӄыльын пэлянэн вэлвынн.
Кыеквъи вэлвын, ӄулильыръуиʼ:
– Кок-кок, эʼми пипиӄылгын?
Ынӄо-ым риʼ'эиʼ вэлвын вээмык гыргоча. 
Рэӈамъянма нинэгитэӄин мимыл. 
Льунин чиниткин выйилвыйил мимлычыку. 
Ӄулилыръуиʼ:
– Ынръам мэӈин? Китак+ун мыйъон!
Йъонэн чиниткин выйилвыйил. 
Аʼйӈавъевыӈонэн чиниткин выйилвыйил:
– Мэй, ӄыетги! Ӄынвэр мэчелкылнин:
– Ынръам мэлгымнин выйилвыйил! Ӄынвэр тэӈэлкылнин. 
Ӄулилыръуиʼ:
– Вынэ, ӄэйвэ гымнин выйилвыйил! Чемэт ынӄэната пипиӄылгын гынтэквъи льукэлиткыльуйгым эʼӄэлиӈу эмлыӈэ!
Ф. Тэӈэтэгын, Чавчывэн лымӈылтэ
