Дина КЭУКЭЙ, авынбиблиограф анадыркэн Публичныкэн библиотекэн нынныльын Тан-Богоразын
Павел Виноградов – тэленъеп гэнъэтлин ыʼлгытумгу морыггазетагты.
Калевэтгавыльа этаны лыги нэлгыркын, иӈӄун газетак нымкыче ынан гатвылен чиниткин космосляйвыгыргын ынкъам ынкэкинэт вагыргыт игыркинэт ынкъам ӈотӄокэнат тэнмычьыт космонавтикэн.
Аймавыӈӈок ынин оʼратъылёӈэт моргынан ытлён мыттэнӄитпыӈыркын ынкъам мытынкэтъоӈатыркын калевэтгавыльэты ынин эргыпатыльын вагыргыръэт.
Павел Виноградов гъурэтлин Магаданык ройыръык инженерэн.
Гэмэйӈэтлин Чукоткак, миӈкы 1970 гивик гэкэлиткуплыткулин Анадыркэн мынгытгэвэкалеткорак №1.
Гэкэлиткулин Москвакэн авиационныкэн институтык факультетык «Летатыльные аппараты».
Ачгыта калеткома ытлён гэмигчирэтлин студентэн конструкторкэн бюрок «Искра», гитлин авынлаборанто ӄол лабораторияк.
Кэлиткуплыткук нанпэлявын институтык рымагтэты мигчирэтык.
Апрелтагнэпы 1977 гивикин Павел Виноградов гамэгчерымголен отраслякэн лабораторияк инженеро ынкъам авнинженеро.
Августык 1983 гивик гамэгчерымголен Ракетныкэн-космическыкэн корпорацияк «Энергия».
Ынан гыму нинэлгыӄин гыюлетык мигчитти ыʼтвыръин «Союз» ынкъам орбитальныкэн ыʼтвин «Буран», лымӈэ ӄутти вагыргыт космосляйвыкэн.
1987 гивик Павел Виноградов гэнъэтлдин отрядык космонавтыргэн, ынан гатаӈынкалыровленат гыёлятгыргыт нъэлкин отрядык, августык-ым 1988 гивик гарылгылен оʼрамръальо итык космонавто.
13 майык 1992 гивик гэнъэтлин кандидато космонавто иткин.
Ӈирэӄ гивиткуӈит гатэнмавлен Центрык тэнмавкэн космонвавтыт.
5 августык 1997 гивик Павел Виноградов Анатолий Соловьёвына рээн гэриӈэлин космосэты ыʼтвэ «Союз ТМ-26».
10 апрелык пытлиӈычьэтыльын космосык лейвык 198 ныкэрэтъылёӈэт Павел Владимирович Виноградов гинэнпиривлин Золотокэн медаля Героен Россиякэн Федерациен.
Мартатагнэпы 1999 гивикин итыркын вице-президенто Федерациен космонавтикэн РФ.
Павел Виноградов космосъытвэпы ӈэръамытлынча гантолен. 2014 гэвэтагнэты ымыльэты ынкы гатвален 38 лиӈыткучьывырӈит ынкъам 25 минутти.
Мартак 2013 гивик гэриӈэлин космосъытва «Союз ТМА-08М» командиро ыʼтвин ынкъам космосляйвынвык МКС-35.
Ынӈингивик ытлён ынанынпычьо космонавто гэнъэтлин – 59 элеӈитыльу.
24 апрелык 2008 гивик гэнинэнпиривлин ордена «За заслуги перед Отечеством  V степени», 22 октябрык 2015 гивик - ордена Мужества.
Рывэтгаквыргыгъет Советэн депутатэн городкэн округэн Анадырь 26 декабрык 2006 гивик Павел Владимирович Виноградов ганэргыпныннатлен Эргыпатыльо гражданино городэн Анадырь.
Космосляйвыма ынан гэнлейвылинэт флаг-кыргычьын Чукоткакэн автономныкэн округэн, газета «Крайний Север» ынкъам чукоткакэн пеликен.
Космосляйвыма ытлён космосъытвэпы гавэтгавлен ӈиныльык рээн.
