Гантэнмавлен Эвын ЭКУКЭКИНЭ
Перевод Амалваӈ вальыт яанаӈат гантомгавленат о´равэтльарык, танляйвыӈ йыркъылгыпы уттынутэк ынкъам эмнуӈкы льэлеӈкы.
Эргыпатыльа учёныйына, этнографа Владилен Леонтьевына, гыютльэ лыгъоравэтльэн-айванальэн культурак ӄол ынин тайкыё кэлиӄэйык «Самый сильный, самый ловкий» гэкэлилин, иӈӄун лыгъоравэтльата ынкъам айванальа нэтэйкынэт вэлвыегыт.
Нытвыӈӈоӄэнат ынӄэнат яанаӈат ӄутырык ракеткано теннисыткукин.
Тайкыёно вэлвыегыт ныяаӄэнат нъумӄинэт вырвыртэ ёмромкэн.
Ынӄэнат нычвиӄинэт гаттэта, ныкылтыӄинэт чьомыткынтэ ынкъам вытгыр кылтыёк нынъылиӄинэт укттытъулти.
Нытомгатӄэн ягпэрагты вальын, кылтэ- ты вальын оттыяанаӈ.
Ынӄоры о´мрынэлга нынтомгавӄэн о´птыма укопрапэральын яанаӈ.
Ынкы ныйпатӄэн гыткалгын лыгъоравэтльэн вэлвыегыткульин.
Вэлвыегыт ралетяанан люӈылгыльыт, ӄаарамка нытэйкыӄинэт тигыт.
Вэлвыегыт ынӈатал плепы вальыт чейвык эмнуӈкы ы´лванвык, аӈӄагыннэгӈыттыльа ынӄэнат таӈъъяаӈ – этэӈӄитыкыльин мэмлыткынгыпы так.
Ыныкит-ым охотник миӈкы ӈан и´рыльылӄыл, вэлвыегыт тэвэнаӈо инэ- эру гитэ.
Пастухо энма гымнан ӄол нинэнтигым нинэнлейвигым ӈалвыльэты рэвылӄэвма, уӈэлык орвъаманма, увиркиплыткук орвыткын нинэтинэӈэгим чывэё уттэ ынкъам нинъэмэтигым ярагты.
