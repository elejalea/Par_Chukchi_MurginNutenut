Эвын ЭКУКЭКИ
Чавчыва рывэнавъё ӈэлвыл  валёмыӈ нынъэлӄин ынкъам ымы гынкыӈ вальо нитӄин.
Бригадир ӄорагынрэтыльэн совхозэʼн нынныльын XXII съездэн КПСС Качьагыргын 1970-ӄавкэнат гивиткук нивӄин: «Этъопэл турэлеръук вэты гыму гэлгэ таӈалвыльыӈгыргын».
Ынӄэн таӈчечавыӈ:  элек торывтатык  ӄаат лымынкыри гарамананчера.
Гырокы  ӄэюут виин  аромкэгты  вальо люӈитэ, гэвиитэ ытльак ӄача.
Омавык-ым ынкъам рораръок гамгота капчачляйвык, гатымӈэва ынкъам гамгота ытльаэнарэрык, эʼмитлёнат (рэквытти) нэмыӄэй гэрынгытвитэ.
Ӈэлвыл ынӄэната ымыльэты гэгынрытвитэ  нэмыӄэй.
Ынӄэн нъэлык чавчыва энмэч тайкыёлӄыл ӈэлвыл.  Ыргынан гатата ӈэлвыл ӄойвэгыргэты, миӈкы эгыӈ гатвата ывнкъам танрылгатык паӈъэвӈытонво.
Ынӈэӈӄач ӈэлвыл гэгынритэ амрытэнма ӈроӄ ныкэрэтъылёӈэт, ванжэван агтатка ӄолеавээнвэты.
Ӈэлвыл вэты ыннанванвык гэгынритэ, иӈкʼун ныкэвыркын чаакайытвак.
«Ынӈэнъылёткок этъопэл авнагтыӈаёвка рытъёлӄыл, вэты чеэкэй вальылӄыл, « - гивалин Качьагыргын.
Виталий Задорин, Гыёлятгыргын Качьагыргынэн, Магаданкэн такнигаӈынвын, 1976 гивиӈит
