Иван О’МРУВЪЕ
О’ткэн гатваленат ытръэч 42 элен’итти, титэ ытлён пэлк’этгъи, э’квыргъам панэна натан’кэтъоркын чукоткальа.
ЭВЫН К’УТТИ К’ОРАГЫНРЭТЫЛЬЫЛК’ЫЛТЭ
1933 гивик О’ткэ, микынэ гэплыткулинэт курсыт вэтгавъёлгыткокэн, гэвинрэтлин рыегтэлевык челюскиныльыт, микынти гэмпэлинэт гэлыткынэты эрэрыльын пароходгыпы, 144 милмил урэльу э’н’ыткынгыпы Увэлен.
Нымкыче ытлён гателеграмматколен вэтгавъёлгэпы гэлыткынкэн лагерэты ынкъам ынк’оры Майн’ынотагты ынк’энат гэнн’ивэ.
Лымн’э ынан гэплыткулинэт курсыт тылечьыткукин рывантыё Чукоткакэн культбазак вальын К’ытрык ынкъам гитлин тылечьыткульу ныппылюк’ин шхунак.
Чама гэмигчирэтлин вэлыткорак’айык, ывинтэтыльу гитлин калеткорак.
Элек охотама нывинрэтк’ин ытлыгэты ан’к’агыннэгн’ыттык.
Пэтле О’ткэ гэнн’ивылин тайкынво вэтгавъёлгыткостанция Ватыркагты, мин’кы нантомгавын Вилюн’эйкин культбаза.
Лейвыльын Ватыркагты О’ткэ ынн’ингивиткук гымнин чычеткин нымнымэты гатвылен ынтуулпырэ А’ляна, микынэ гаматален гымнин чакыгэт Люба.
Алексей Павловичын галяльын гивик гэнъэтлинэт 94 элен’итти, вачак’ панэна ынан игыр лыги лын’ыркынин етыльын Ватыркагты О’ткэ.
А’ля нивк’ин, энмэн ытлён н’ирэче гэгынтэвлин интернатгыпы амнон’эты н’алвыльэты эмъэнк’этык кэлиткук.
О’ткэна, лыги лын’кы ынк’эн, кэлиныгйивэтыльыт ивнинэт, опопы мачынан А’ля эвнэнкэлиткувкэ, к’элюк’ эвын к’утти мэйн’этыльылк’ылти к’орагынрэтыльо.
ЭНМА ЫТЛЁН ПРЕДСЕДАТЕЛЁ
Чинит гымнан О’ткэ эльукыльин.
Э’квыргъам лыги гымнан ымыльо ынинэт н’ээккэт.
Энмэчевын к’ол ынин н’ээккэк – Надяна рээн 60-к’авкэнат гивиткук гэкэлиткуйгым Анадыркэн педучилищек Айгыск’ываратыргэн ынкъам нымкыче гавалёмлен тывъё ынин ытлыгын каленыгъеватыльэпы ынкъам ынпыянвэпы.
Н’ээккэт О’ткэн гэмэйн’инъэтэтлинэт мэйн’этык.
Ынн’ин, Надежда О’ткэ 1980-1990 гивиткун’ит гитлин председателё Чукоткакэн окрисполкомэн, гэнъэтлин кандидато историческыкэн наукэн.
К’утти вагыргыт О’ткэн гымнан гэйгулетлинэт ынпыянвэпы ынкъам ынин н’авъангыпы – Лемма Магометовнайпы.
Гымнан к’улин нинэльуйгым н’аргын вальын ченэтрак к’ача Лемма Магометовна.
Нэймэвигым ыныкы ынкъам нымгоморэ пычвэтгавык лыгъоравэтльелымэл – Лемма Магометовнана, айванальын’ава, гэтэн’ыйгулетлин лыгъоравэтльэн йилыйил.
Нымытвавагыргын О’ткэн гэкэлилин нымк’ыкин кэлик.
Вэнлыги-ым, антыяаткэгты, чымк’ык мытвыгъан.
1946 гивик нымытвальа нымнымкин Эк’к’эни О’ткэ гэльулин депутато Верховныкэн Советэн СССР Чукоткакэн национальныкэн округгыпы.
Ытлён ынкы гэмигчирэтлин 1946 гэвэтагнэпы 1954 гэвэтагнэты.
1947 гивик О’ткэ гэнъэтлин председателё Чукоткакэн округкэн исполкомэн.
Ытлён гинъэтэтлин раройвавынво экономика Чукоткакэн: мэгчерымгогъат нотагаймычьыэнарэркэнат партият льонво золото; гантомгавлен Чукоткакэн таран’управление, раройвавынво пылвынтынтокэн промышленность гатайкымголенат посёлок Эквыкыннот, ымыск’ыльын ан’к’аы’тымпан; гэнмэйн’эвлинэт ан’к’аы’тымпанвыт Провиденияк, Пээкик, Бухтак Угольная.
О’ткэ гаванлялен Советкэн правительствогты рытомгавынво округык подразделение Гражданкэн авиациен.
1947 гэвэтагнэпы моогъат рин’элейвык округык ынкъам Хабаровскэты, Магаданэты ынкъам Москвагты.
Сельскакэн хозяйствок аройвавымгогъэ тан’алвыльын’гыргын к’орагынрэтынвык, мыкатымгогъат ан’к’агыннэгн’ыттыкэнат колхозтэ, тэннын’кинэт артельтэ.
Колхозникыльэты Чукоткагты наныпкэратын’н’онат рымыльава рытыльыт нымытварак’агтэ; ан’к’агыннэгн’ыттыльэты нэныпкирэтынэт торвельботтэ, нымкык’ин нымнымыткук мэгчерымгогъат зверофермат; Анадыркэн районык намгонат рынн’эвык роолк’ыловощит.
Мигчир О’ткэн энма председателё окрисполкомэн ганъялен Правительствота – декабрык 1950 гивик ытлён гинэнпиривлин ордена Ленинын.
Справка «КС»
Июлык 1947 гивик исполком Анадыркэн Советэн депутатыргэн мэгчетльываратэн гавэтгыльатлен: «Тан’кэтъонво чит итыльын председателё Чукоткакэн окрисполкомэн О’ткэ равытгыр Строительная – ныннэтык равытгыро О’ткэн».
