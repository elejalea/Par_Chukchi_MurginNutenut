Ирина РОМАНОВА, заместитель директорэн Музейныкэн Центрэн «Наследие Чукотки»
Перевод Кэлиткуплыткульын историческыкэн факультетык Ленинградкэн университетэн, энмэч гыютльэн нотагаймычьыэнарэрынвык мигчирэтык Арменияк, Туркменистанык, Забайкальек, кандидат историческыкэн наукэн, э´квыргъам еп нылгиныӈинӄин ытлён 1955 гивик гамэгчерымголен тэӈытръэчкин ынӈингивик музейык Чукоткакэн национальныкэн округкэн Мытлыӈэн гивиӈит ынкэкинэт яанаӈт ӈирэче мыкыӈ гэтчылинэт.
ЯРАӇЫ, МИӇКЫ ТАНЛЬОӇ ИМЫРЪЭНУТ
Кэлик ынан тайкыёк «По следам древних костров» гатвылен музей 1950-ӄавкэнат гивиткукин ынкъам гэныгйивэтлинэт мигчитлыӄылти ынӄэн раройвавынво, рымкавынво ынкэкинэт яанаӈат таляӈкэнавагыргыкэнат.
Ынан гэкэлилин: «Чукоткак варкын музей, яраӈы, миӈкы, нивӄинэт лыгъоравэтльат, танльоӈ имыръэнут, яаё ы´ттъытльэ тэлеӈкы.
Ынӄэн яраӈы гэтэйкылин ромотта 1930-ӄавкэнат гивиткук ынкъам чьувылтэтыркын мыкэтык яанаӈат ромакавъёттэ.
Энмэч ӈыраӄ гивиткуӈит музея рылеркынинэт археологическыкэн ноталяйвыгыргыт, ӄымэл-ым мытыйгулетыркынэт тэлеӈкинэт вагыргыт авыннымытвальэн ӈутиннутэк» – гэкэлилин Николай Диковына.
Диков мэгчеранма музейык ныкытрэватӄэн.
Ынӈин, 1956-1959 гивиткуӈит ынан моонэнат гыюлетык нутэйиквит Чукоткакэн, аӈӄачормыкэнат нымытваванвыт ы´ттъыютльин, гыюленнинэт ваамъёчгыт Анадырэн, О´мваамэн, Ваӈӄарэмакэн, льунинэт нымытваванвыт ы´ттъыютльин гытгык ӄача Красное ынкъам Чировое.
Ынан льунинэт нымкыӄин панэнаванвыт тэлеӈкинэльин, титэ ынӄэнат гатваленат.
Ынан гэкэлилин, иӈӄун культура лыгъоравэтльаваратэн ынкъам аӈӄагыннэгӈыттыльэн ынкъам ынныӈыттыльин эвын гатвален II-I векык унмытэленъеп, миӈкы ынанъыттъыёл нымытвальо гитлинэт янор лыгъоравэтльэн ы´ттъыютльэт.
Рыйголявъё антрополога-учёныя М. М. Герасимовына – Г. В. Лебединскаяна лявтыы´тъымгыпы гэныгйивэтлин вальын льулӄыл ынкъам игыр танльоӈ ынӄэн Аналддыркэн музейык миӈкри вальо гатвален о´равэтльан ӈроӄ тысячтэ гивиӈитти яалегты.
ЯАНАӇАТ – ЭВЫНКУМЪЫН МУЗЕЕН
Диковына лымӈэ гамголен гыюлетык тэлеӈкин айванальэн культура.
1969 гивик ынан гэльулин ӄытрыкин панэнаванвык аӈӄальэн яаё ваӈӄытъяанаӈ гыннигӈыттыкин.
Диков гивлин, иӈӄун культура тэлеӈкин аӈӄагыннэгӈыттыльэн микынэ люнрэтыльын Чукоткагты, ипэ ынӄэн гатомгатлен Эйгысӄык.
1956–1959 гивиткуӈит гэнумэкэвлинэт льоёттэ нымкыӄин тэлеӈкы яаёттэ яанаӈат.
Ынӈингивиткуӈит гэльулинэт мыкыӈ 1.5 тысячкэнак яанаӈат.
Лымӈэ игыр музейык варкыт нымкыӄин виилыгтыт, тайкыёттэ вама ынӄэнат ноталяйвыгыргыт мигчитльин музейкин.
Николай Диков эмэлкэ итыркын ы´ттъыёлкэн директоро округкэн музеейык, микынэ ромакавымгонэнат льоёттэ яанаӈат тэлеӈкинэт ынкъам ынӄэнат тывнэнат наукгъет.
Ынан гэнӄитпэвлинэт винрэтык ытлён румэвык яанаӈат тэлеӈкинэт эвынӈуткэкинэт нымытвальыт.
Гамгаляйвынвэпы ынан тэӈэвын нинэрэтӄинэт ынӄэнат ынкъам нэнамгоӄэнат гыюлетык.
Мытлыӈэн гивиткуӈит мигчирэткин директоро музейык ынкы гатваӈӈоленат ӈирэче мыкыӈ яанаӈат льоёттэ.
Учёныен, гыютльин тэлеӈкинэт культурак ынкъам археологияк Северо-Востокэн Россиен, членэн-корреспондентэн Россиякэн академиен наукэн, профессорэн Николай Николаевич Диковын (1925–1996) 17 мартак нъынъэлынэт 95 гивиӈитти о´раттагнэпы.
ПАГЧЕӇГЫРГЫТ ТАЛЯӇКЭНАВАГЫРГЫТ
Энмэч мэгчеранма Магаданык Николай Диков гатвален икутъэр ноталяйвынвык гыёлятынво тэлеӈкинэт вагыргыт авынчукоткальэн.
Нотаргыткогыргыт ынан гэнлелинэт ваамъёчгык Анадырваамэн, О´мваамэн, Пенжинан ынкъам ы´ттъыютльин айванальэн Увэлек ӄача, Чиник, Чегтук ӄача 1960-ӄавкэнат гивиткук.
1967–1968 гивиткук Николай Никлаевичына гыёлятымгонэнат энмыкэнат рисугнкат ынкъам ӈирэӄ унмытэлеӈкинэт ралӄаӈынвыт Эйгысӄык.
Ынан гэльулинэт мыкыӈ мытлыӈӄлеккэнак рисункат, тайкыёттэ энмык тэлеӈкинэт гыннигӈыттыльэ.
Ымыльо льоёттэ энмык Диковына гатвыленат кэлик, тайкыё 1971 гивик «Наскальные загадки древней Чукотки».
Ынӄэнат энмыкэнат рисункат ымы игыр пэгчиӈу нэлгыркынэт учёныйрык ынкъам э´йӈэвыткуркыт ырыкы вак ынӈэнӄач нутэлейвык таӈыйголятынво тэлеӈинэт вагыргыт эвынӈуткэкыльин.
Лымӈэ ӄол ляйвыгыргын гатвален Диковын 1975 гивик Омӄэлерэты, титэ мачалваӈ гэвытрэтлин таляӈкэнавагыргын айванальэн.
Ынӄэн ляйвынвык гатвален ынин гыюлетыльын Тэйр Тасян.
Эмӄитпыльэтык ынкъам инъэтэтк Николай Диков Чукоткакэн округкэн музея моонэнат тэйык чиниткинэт «Записки…».
Ынӄэн, этъыманы, тэӈытрэчкин ынӈингивик Чукоткак наукагъёляткэн кэликэл-журнал.
Николай Николаевичына гэнӄитпэвлинэт ӄутти о´равэтльат нэмыӄэй гыюлетык таляӈкэнавагыргыт Чукоткак.
Тэнмычьо, Маргарита Александровна Кирьяк мигчитльэрык рээн музейкин гатваленат О´мваамык ынкъам гытгык Эӄитыки, миӈкы гэльулинэт лымӈэ ӄутти тэлеӈкинэт яанаӈат эвынӈуткэкыльин.
Нынны Николай Николаевичын эргыпатэты натвыркын яатльа Чукоткакэн, миӈкрик ӄун ынан гэйгулетлинэт нымкыӄин вагыргыт вальыт ы´ттъытльин.
Редакторо итык ытлён 1989 гивик гэтэйкылин кэликэл «История Чукотки с древнейших времён до наших дней».
