Эвын ЭКУКЭКИ
Перевод Кэлик «Ынӈин гатвален…» Тасян Теинына гатвылен таройыръыӈгыргын айванальэн тэлеӈкы.
Ройыръык айванальэн гатвата ы’вэӄуч, ӈэвъэн ынкъам кмиӈыт.
Ыныкит яраӈы ныркывӄэн, ырыгрээн ганымытвата ынпэвыльыт йытоткольыт.
Ыныкит пэлӄэтыльыт йытоткольыт гитлинэт чычеткинэльу, пэлятыльыт ейвэлти нынъэлӄинэт йичьэмиттумгу ынкъам чакэттомго кмэӈэты ройыръэн.
Ынӄэнат кмиӈыт айванальа нытвыӄэнат анлисаг’аӄ.
Кмэӈынмайӈаквыргын ейвэлык гамыкытвален Аляскальык.
Гаймычьыройыръык, миӈкы авынральын нитӄин кынтэгыннигӈыттыльу, ӄол гитэ ӄляволен гатвата ӈирэют лымэвыр мыкыӈ ӈэвъэнти.
Ынпычьын ӈэвъэн нитӄин авынэтынво ярамэгчерык.
Ынан нинэнмэйӈэвӄинэт чиниткинэт ынкъам ӈинчьин кмиӈыт.
Ӈинчьэт ӈэвъэнти нываӈэӄэнат, нывиӄинэт, нытэнэлгыӈӄинэт, нинээнӈэтӄинэт тымъёк гынникык.
Ӈэвъэнти натчьатӄэнат ыннэн ёрочыко, э’квыргъам ымыльо рыгъеватъё чиниткин ванвык.
Ӈинчьэн ӈэвъэн вэты ӄырымэн а’рэткочьо итыльылӄыл мигчирык ынпычьин ӈэвъэнин.
Ыныкит ы’ттъыёлкэн ӈэвъэн уйӈэ экмиӈыкэ гатвален, ӄлявол гаймаӈэн лымӈэ гэӈирэӄэвэ ӈавтыӈык.Тэнмычьо, ы’ттъыёлкэн илирык нымытвамгольэн Таянын гатваленат ӈирэӄ ӈэвъэнти.
Ӄлявол ‘ырымэн ярамэгчерык рэӄыльылӄыл, ӈэвысӄэт-ым ӄырымэн гыннигӈыттыльу итыльылӄыл, ынӄэн амӄляволен мгчир.
Ынӈин тымӈалголяӄ ринӈыльыт ӄлявол лымэвыр ӈэвысӄэт чычеткинэльу ивыну гэлгэ ынкъам э’ӄэлтэтыльу ройыръывагыргык.
Лыгэн-ым, ӈиныльин ӈэвъэнин гатваленат нымкыӄин мигчитти ратвакэн.
А’нӄатгыргын ройыръытвак нырылгыӄэн тэнанъаӄаӈгырго ройыръытвагыргык.
Ӈинчьэт ӈэвъэнти а’ӄантыӈ ройыръэпы.
Ынинэт кмӈыт ӄынвэр гэкэвэ мэйӈэтык ынпычьыӈэвъэнык, микынэ ытри гэнмэйӈэвэ.
