1982 гивик Магаданкэн такнигаӈынвык гэтэйкылин кэликэл гастихма дальневостоккэн поэтэн Владимир Першинын, миӈкы ынан вэтгаво гэлгылин ы’лгыльатгыргын - О’ратнотагты , Айгысӄынотагты, э*митлён ынык гитлин ӄэтпыкво нымытвак, ытлыгыргин ванвэты, ытльагты, ӈавысӄатэты – лыгэн-ым ымыльорыкы ынкъам эмыраӄэты.
Ынӄэн кэлик гайпатленат ымы стихыт елыльатъёттэ тэкэлиӈыльэ лыгъоравэтльэн поэтыргэн, ымы Клавдия Гэутваалын, микын ӄол стихотворение мыткалейпатыркын.
