Дина КЭУКЭЙ, Иван О´МРУВЪЕ
Перевод Энмэч 31 гивиӈитти анадыркэн Публичныкэн библиотека итыркын нынныльу Владимир Германович Тан-Богоразын, ынин о´ратъылёӈэттагнэпы 27 апрелык галягъат 155 гивиӈитти, Еп январык ӈутингивикин ынкы гэтэйкылин выставка, рыгъевавынво ынӄэн таӈэргыпатыльын о´равэтльан, мэӈин гинъэтэтлин рымагтэты раройвавык культура ынкъам таӈвагыргыт айгысӄываратыргэн Россиен.
Ынӄэн выставка ратвагъа ымыльэты ӈотӄэн гивиӈит.
Вальын студентэн вэчыёгты а´рӄачьатгыргык Богораз рытымучьэвэ гэпирилин ынкъам гавосӄырален янор Петропавловскыкэн крепостык, 1886 гивик-ым гэнэквэтэвлин танымчаӈынво Средне-Колымскэты.
Вама ынкэкин нутэк Богоразына моонэнат гыюлетык нымытвавагыргыт, ынӈатал энъататэты, рыпэтым 1894 гивик ытлён нэмыӄэй 7 натвыгъан этыльу эноталяйвынвэты гыёлятынво вагыргыт лыгъоравэтльэн ынкъам ӄутти варатыргэн Северо-Востокэн Евразиен.
12 тысячтэ вёрстыт яанэнат Богоразына ӈирэӄ гачывэптыма гивиӈит ноталяйвыма Экулымэк ынкъам Чукоткак.
Льоёттэ вагыргыт ынан ӈотӄоры гэкэлилинэт рассказык.
Ынан гыюленнинэт лыгъоравэтльэн ынкъам айванальэн йилыт.
Э´квыргъам ытлён гатаӈэргыпатлен титэ тэйкынин мэйӈыкэликэл «Чукчи», миӈкы гатваленат ӈроӄ разделтэ – «Социальная организация», «Религия» ынкъам «Материальная культура» нымкъэв гатвылен нымытвавагыргын эвынӈуткэкыльин талпытыляма XIX век ынкъам энэнэма XX век.
Наӄам варкыт тайкыёттэ виилыгтыт, ымы лыгъорапвэтльак рээн ноталяйвыама.
Ы´ттъыёлкэн разделык Владимир Германович Тан-Богоразына гатвыленат, миӈкы нымытваркыт ынкэкинэт о´равэтльат, миӈкыри вальыт ытри, о´ратгыргыт ыргинэт, ӈавтыӈгыргын ыргин, ройыръыт, правот ыргинэт.
Ынӄэн раздел гэтэйкылин янор англияльэн йилымил Нью-Йиоркык 1904–1909 гивиткук, русильымил – Ленинградык 1934 гивик.
Ӈирэӄэв раздел «Религия» янор гэтэйкылин англияльэн йилымил 1912 гивик, русильин йилымил – 1939 гивик.
Ынӄэн разделык гатвыленат кальатаароӈгыргыт, гыргыртэ, нымкъэв гатвыленат крычмыт, аӈаӈыткогыргыт эмыръатаароӈгыргыт авыннымытывальэн ынӈиннутэк, о´ратгыргыт ынкъам уйӈэ нъалгыргыт о´равэтльэн .
Разделык «Материальная культура» гатвыленат ӄорагынрэтгыргын, таы´ттыӈгыргын, гыннэгӈыттыгыргын ынкъам ынныӈыттыгыргын.
Лымӈэ миӈкри вальыт лыгъоравэтльэн нымытварат, яраяанаӈат, роолӄылтэ, мигчир, эвиръыт, увичвыт, крычмыт.
Чиниткинэт пыӈылтэлык Владимир Тан-Богоразына гатвыленат нымытвавагыргыт .
Ынин монография «Чукчи» эргыпатыркын ынкъам Владимир Германович Тан-Богораз итыркын ӄол гыютльу этнографо ымнотаеквэкэн учёныйырык.
Ытлён гэпэлӄэтлин 1936 гивик.
Гэнумкэвлин Ленинградык.
Лымӈэ
Таӈыйголятынво культура ынкъам вагыргыт эвынӈуткэкыльин, калейпатъёттэ монографияк «Чукчи», романык «Восемь племён», «Союз молодых», «Жертвы дракона», пыӈылтэлык «Мёртвое стойбище», «Кривоногий» ынкъам ӄутти, тэкэлиӈыльэ ӈотӄэн статьяк ӄол гэнтэ гапытӄыкалевэтгава Тан-Богораз.
